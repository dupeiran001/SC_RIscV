module pc(
  input         clock,
  input         reset,
  input  [7:0]  io_pc_ctrl,
  input  [31:0] io_pc_imm,
  output [31:0] io_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc_reg; // @[pc.scala 17:19]
  reg  tmp; // @[pc.scala 18:16]
  wire  _T_2 = 8'h0 == io_pc_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _pc_reg_T_1 = pc_reg + 32'h4; // @[pc.scala 29:24]
  wire  _T_3 = 8'h3 == io_pc_ctrl; // @[Conditional.scala 37:30]
  wire  _T_4 = 8'h1 == io_pc_ctrl; // @[Conditional.scala 37:30]
  wire  _T_5 = 8'h2 == io_pc_ctrl; // @[Conditional.scala 37:30]
  wire  _T_6 = 8'h4 == io_pc_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_0 = _T_6 ? io_pc_imm : pc_reg; // @[Conditional.scala 39:67 pc.scala 41:14 pc.scala 17:19]
  wire [31:0] _GEN_1 = _T_5 ? io_pc_imm : _GEN_0; // @[Conditional.scala 39:67 pc.scala 38:14]
  wire [31:0] _GEN_2 = _T_4 ? io_pc_imm : _GEN_1; // @[Conditional.scala 39:67 pc.scala 35:14]
  wire  _GEN_5 = ~tmp | tmp; // @[pc.scala 24:26 pc.scala 25:9 pc.scala 18:16]
  assign io_pc = pc_reg; // @[pc.scala 20:9]
  always @(posedge clock) begin
    if (reset) begin // @[pc.scala 21:21]
      pc_reg <= 32'h0; // @[pc.scala 22:12]
    end else if (!(~tmp)) begin // @[pc.scala 24:26]
      if (_T_2) begin // @[Conditional.scala 40:58]
        pc_reg <= _pc_reg_T_1; // @[pc.scala 29:14]
      end else if (_T_3) begin // @[Conditional.scala 39:67]
        pc_reg <= io_pc_imm; // @[pc.scala 32:14]
      end else begin
        pc_reg <= _GEN_2;
      end
    end
    if (reset) begin // @[pc.scala 21:21]
      tmp <= 1'h0; // @[pc.scala 23:9]
    end else begin
      tmp <= _GEN_5;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  tmp = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module alu(
  input  [7:0]  io_alu_ctrl,
  input  [31:0] io_alu_src_1,
  input  [31:0] io_alu_src_2,
  output [31:0] io_alu_out
);
  wire  _T = 8'h0 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _io_alu_out_T_1 = io_alu_src_1 + io_alu_src_2; // @[alu.scala 20:34]
  wire  _T_1 = 8'h6 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _io_alu_out_T_2 = io_alu_src_1 & io_alu_src_2; // @[alu.scala 23:34]
  wire  _T_2 = 8'h1 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _io_alu_out_T_4 = io_alu_src_1 - io_alu_src_2; // @[alu.scala 26:34]
  wire  _T_3 = 8'h5 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _io_alu_out_T_5 = io_alu_src_1 | io_alu_src_2; // @[alu.scala 29:34]
  wire  _T_4 = 8'h7 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire [94:0] _GEN_26 = {{63'd0}, io_alu_src_1}; // @[alu.scala 32:34]
  wire [94:0] _io_alu_out_T_7 = _GEN_26 << io_alu_src_2[5:0]; // @[alu.scala 32:34]
  wire  _T_5 = 8'h8 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _io_alu_out_T_9 = io_alu_src_1 >> io_alu_src_2[5:0]; // @[alu.scala 35:34]
  wire  _T_6 = 8'h9 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _io_alu_out_T_13 = $signed(io_alu_src_1) >>> io_alu_src_2[5:0]; // @[alu.scala 38:73]
  wire  _T_7 = 8'h4 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _io_alu_out_T_14 = io_alu_src_1 ^ io_alu_src_2; // @[alu.scala 41:34]
  wire  _T_8 = 8'h2 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire  _T_11 = $signed(io_alu_src_1) < $signed(io_alu_src_2); // @[alu.scala 44:34]
  wire  _T_12 = io_alu_src_1 > io_alu_src_2; // @[alu.scala 47:25]
  wire  _GEN_1 = io_alu_src_1 > io_alu_src_2 ? 1'h0 : _T_11; // @[alu.scala 47:40 alu.scala 48:20]
  wire  _T_13 = 8'h3 == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire  _T_14 = io_alu_src_1 < io_alu_src_2; // @[alu.scala 52:25]
  wire  _GEN_3 = _T_12 ? 1'h0 : _T_14; // @[alu.scala 55:40 alu.scala 56:20]
  wire  _T_16 = 8'ha == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire  _T_17 = io_alu_src_1 == io_alu_src_2; // @[alu.scala 61:25]
  wire  _T_18 = 8'hc == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire  _T_19 = io_alu_src_1 != io_alu_src_2; // @[alu.scala 68:25]
  wire  _T_20 = 8'hd == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire  _T_24 = 8'hb == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire  _T_27 = $signed(io_alu_src_1) >= $signed(io_alu_src_2); // @[alu.scala 82:34]
  wire  _T_28 = 8'he == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire  _T_30 = 8'hf == io_alu_ctrl; // @[Conditional.scala 37:30]
  wire  _T_31 = io_alu_src_1 >= io_alu_src_2; // @[alu.scala 96:25]
  wire  _GEN_10 = _T_30 & _T_31; // @[Conditional.scala 39:67 alu.scala 16:14]
  wire  _GEN_11 = _T_28 ? _T_14 : _GEN_10; // @[Conditional.scala 39:67]
  wire  _GEN_12 = _T_24 ? _T_27 : _GEN_11; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_20 ? _T_11 : _GEN_12; // @[Conditional.scala 39:67]
  wire  _GEN_14 = _T_18 ? _T_19 : _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_15 = _T_16 ? _T_17 : _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_16 = _T_13 ? _GEN_3 : _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_17 = _T_8 ? _GEN_1 : _GEN_16; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_18 = _T_7 ? _io_alu_out_T_14 : {{31'd0}, _GEN_17}; // @[Conditional.scala 39:67 alu.scala 41:18]
  wire [31:0] _GEN_19 = _T_6 ? _io_alu_out_T_13 : _GEN_18; // @[Conditional.scala 39:67 alu.scala 38:18]
  wire [31:0] _GEN_20 = _T_5 ? _io_alu_out_T_9 : _GEN_19; // @[Conditional.scala 39:67 alu.scala 35:18]
  wire [94:0] _GEN_21 = _T_4 ? _io_alu_out_T_7 : {{63'd0}, _GEN_20}; // @[Conditional.scala 39:67 alu.scala 32:18]
  wire [94:0] _GEN_22 = _T_3 ? {{63'd0}, _io_alu_out_T_5} : _GEN_21; // @[Conditional.scala 39:67 alu.scala 29:18]
  wire [94:0] _GEN_23 = _T_2 ? {{63'd0}, _io_alu_out_T_4} : _GEN_22; // @[Conditional.scala 39:67 alu.scala 26:18]
  wire [94:0] _GEN_24 = _T_1 ? {{63'd0}, _io_alu_out_T_2} : _GEN_23; // @[Conditional.scala 39:67 alu.scala 23:18]
  wire [94:0] _GEN_25 = _T ? {{63'd0}, _io_alu_out_T_1} : _GEN_24; // @[Conditional.scala 40:58 alu.scala 20:18]
  assign io_alu_out = _GEN_25[31:0];
endmodule
module ctrl(
  input  [31:0] io_instruction,
  output [7:0]  io_pc_ctrl,
  output [7:0]  io_imm_ctrl,
  output [7:0]  io_data_ctrl,
  output [7:0]  io_select_ctrl,
  output [7:0]  io_reg_ctrl,
  output [7:0]  io_alu_ctrl
);
  wire  _T_1 = 7'h63 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h0 == io_instruction[14:12]; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h5 == io_instruction[14:12]; // @[Conditional.scala 37:30]
  wire  _T_5 = 3'h7 == io_instruction[14:12]; // @[Conditional.scala 37:30]
  wire  _T_6 = 3'h4 == io_instruction[14:12]; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h6 == io_instruction[14:12]; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h1 == io_instruction[14:12]; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_0 = _T_8 ? 4'hc : 4'h0; // @[Conditional.scala 39:67 ctrl.scala 51:23 ctrl.scala 24:15]
  wire [3:0] _GEN_1 = _T_7 ? 4'he : _GEN_0; // @[Conditional.scala 39:67 ctrl.scala 48:23]
  wire [3:0] _GEN_2 = _T_6 ? 4'hd : _GEN_1; // @[Conditional.scala 39:67 ctrl.scala 45:23]
  wire [3:0] _GEN_3 = _T_5 ? 4'hf : _GEN_2; // @[Conditional.scala 39:67 ctrl.scala 42:23]
  wire [3:0] _GEN_4 = _T_4 ? 4'hb : _GEN_3; // @[Conditional.scala 39:67 ctrl.scala 39:23]
  wire [3:0] _GEN_5 = _T_3 ? 4'ha : _GEN_4; // @[Conditional.scala 40:58 ctrl.scala 36:23]
  wire  _T_9 = 7'h13 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h2 == io_instruction[14:12]; // @[Conditional.scala 37:30]
  wire  _T_13 = 3'h3 == io_instruction[14:12]; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_6 = io_instruction[30] ? 4'h9 : 4'h8; // @[ctrl.scala 93:11 ctrl.scala 94:25 ctrl.scala 97:25]
  wire [1:0] _GEN_7 = _T_4 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 ctrl.scala 91:23 ctrl.scala 20:15]
  wire [3:0] _GEN_8 = _T_4 ? _GEN_6 : 4'h0; // @[Conditional.scala 39:67 ctrl.scala 24:15]
  wire [3:0] _GEN_9 = _T_8 ? 4'h7 : _GEN_8; // @[Conditional.scala 39:67 ctrl.scala 87:23]
  wire [1:0] _GEN_10 = _T_8 ? 2'h0 : _GEN_7; // @[Conditional.scala 39:67 ctrl.scala 88:23]
  wire [3:0] _GEN_11 = _T_5 ? 4'h6 : _GEN_9; // @[Conditional.scala 39:67 ctrl.scala 83:23]
  wire [1:0] _GEN_12 = _T_5 ? 2'h0 : _GEN_10; // @[Conditional.scala 39:67 ctrl.scala 84:23]
  wire [3:0] _GEN_13 = _T_7 ? 4'h5 : _GEN_11; // @[Conditional.scala 39:67 ctrl.scala 79:23]
  wire [1:0] _GEN_14 = _T_7 ? 2'h0 : _GEN_12; // @[Conditional.scala 39:67 ctrl.scala 80:23]
  wire [3:0] _GEN_15 = _T_6 ? 4'h4 : _GEN_13; // @[Conditional.scala 39:67 ctrl.scala 75:23]
  wire [1:0] _GEN_16 = _T_6 ? 2'h0 : _GEN_14; // @[Conditional.scala 39:67 ctrl.scala 76:23]
  wire [3:0] _GEN_17 = _T_13 ? 4'h3 : _GEN_15; // @[Conditional.scala 39:67 ctrl.scala 71:23]
  wire [1:0] _GEN_18 = _T_13 ? 2'h0 : _GEN_16; // @[Conditional.scala 39:67 ctrl.scala 72:23]
  wire [3:0] _GEN_19 = _T_12 ? 4'h2 : _GEN_17; // @[Conditional.scala 39:67 ctrl.scala 67:23]
  wire [1:0] _GEN_20 = _T_12 ? 2'h0 : _GEN_18; // @[Conditional.scala 39:67 ctrl.scala 68:23]
  wire [3:0] _GEN_21 = _T_3 ? 4'h0 : _GEN_19; // @[Conditional.scala 40:58 ctrl.scala 63:23]
  wire [1:0] _GEN_22 = _T_3 ? 2'h0 : _GEN_20; // @[Conditional.scala 40:58 ctrl.scala 64:23]
  wire  _T_21 = 7'h67 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire  _T_22 = 7'h3 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_23 = _T_12 ? 3'h5 : 3'h0; // @[Conditional.scala 39:67 ctrl.scala 131:24 ctrl.scala 21:16]
  wire [2:0] _GEN_24 = _T_4 ? 3'h7 : _GEN_23; // @[Conditional.scala 39:67 ctrl.scala 128:24]
  wire [2:0] _GEN_25 = _T_8 ? 3'h4 : _GEN_24; // @[Conditional.scala 39:67 ctrl.scala 125:24]
  wire [2:0] _GEN_26 = _T_6 ? 3'h6 : _GEN_25; // @[Conditional.scala 39:67 ctrl.scala 122:24]
  wire [2:0] _GEN_27 = _T_3 ? 3'h3 : _GEN_26; // @[Conditional.scala 40:58 ctrl.scala 119:24]
  wire  _T_29 = 7'h6f == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire  _T_30 = 7'h33 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_30 = _T_5 ? 3'h6 : 3'h0; // @[Conditional.scala 39:67 ctrl.scala 182:23 ctrl.scala 24:15]
  wire [2:0] _GEN_31 = _T_7 ? 3'h5 : _GEN_30; // @[Conditional.scala 39:67 ctrl.scala 179:23]
  wire [3:0] _GEN_32 = _T_4 ? _GEN_6 : {{1'd0}, _GEN_31}; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_33 = _T_6 ? 4'h4 : _GEN_32; // @[Conditional.scala 39:67 ctrl.scala 168:23]
  wire [3:0] _GEN_34 = _T_13 ? 4'h3 : _GEN_33; // @[Conditional.scala 39:67 ctrl.scala 165:23]
  wire [3:0] _GEN_35 = _T_12 ? 4'h2 : _GEN_34; // @[Conditional.scala 39:67 ctrl.scala 162:23]
  wire [3:0] _GEN_36 = _T_8 ? 4'h7 : _GEN_35; // @[Conditional.scala 39:67 ctrl.scala 159:23]
  wire [3:0] _GEN_37 = _T_3 ? {{3'd0}, io_instruction[30]} : _GEN_36; // @[Conditional.scala 40:58]
  wire  _T_44 = 7'h23 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_38 = _T_12 ? 4'hc : 4'h0; // @[Conditional.scala 39:67 ctrl.scala 200:24 ctrl.scala 21:16]
  wire [3:0] _GEN_39 = _T_8 ? 4'hb : _GEN_38; // @[Conditional.scala 39:67 ctrl.scala 197:24]
  wire [3:0] _GEN_40 = _T_3 ? 4'ha : _GEN_39; // @[Conditional.scala 40:58 ctrl.scala 194:24]
  wire  _T_49 = 7'h17 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire  _T_50 = 7'h37 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_42 = _T_50 ? 4'he : 4'h0; // @[Conditional.scala 39:67 ctrl.scala 214:20 ctrl.scala 21:16]
  wire [3:0] _GEN_43 = _T_50 ? 4'h9 : 4'h0; // @[Conditional.scala 39:67 ctrl.scala 215:19 ctrl.scala 20:15]
  wire [3:0] _GEN_44 = _T_50 ? 4'h8 : 4'h0; // @[Conditional.scala 39:67 ctrl.scala 217:19 ctrl.scala 23:15]
  wire [3:0] _GEN_46 = _T_49 ? 4'hd : _GEN_42; // @[Conditional.scala 39:67 ctrl.scala 206:20]
  wire [3:0] _GEN_47 = _T_49 ? 4'h8 : _GEN_43; // @[Conditional.scala 39:67 ctrl.scala 207:19]
  wire [1:0] _GEN_48 = _T_49 ? 2'h3 : 2'h0; // @[Conditional.scala 39:67 ctrl.scala 208:18]
  wire [3:0] _GEN_49 = _T_49 ? 4'h7 : _GEN_44; // @[Conditional.scala 39:67 ctrl.scala 209:19]
  wire [3:0] _GEN_51 = _T_44 ? 4'h7 : _GEN_47; // @[Conditional.scala 39:67 ctrl.scala 188:19]
  wire [1:0] _GEN_52 = _T_44 ? 2'h0 : _GEN_48; // @[Conditional.scala 39:67 ctrl.scala 189:18]
  wire [3:0] _GEN_53 = _T_44 ? 4'h6 : _GEN_49; // @[Conditional.scala 39:67 ctrl.scala 190:19]
  wire [3:0] _GEN_54 = _T_44 ? _GEN_40 : _GEN_46; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_55 = _T_30 ? 4'h9 : _GEN_54; // @[Conditional.scala 39:67 ctrl.scala 144:20]
  wire [3:0] _GEN_56 = _T_30 ? 4'h6 : _GEN_51; // @[Conditional.scala 39:67 ctrl.scala 145:19]
  wire [1:0] _GEN_57 = _T_30 ? 2'h0 : _GEN_52; // @[Conditional.scala 39:67 ctrl.scala 146:18]
  wire [3:0] _GEN_58 = _T_30 ? 4'h5 : _GEN_53; // @[Conditional.scala 39:67 ctrl.scala 147:19]
  wire [3:0] _GEN_59 = _T_30 ? _GEN_37 : 4'h0; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_60 = _T_29 ? 4'h0 : _GEN_59; // @[Conditional.scala 39:67 ctrl.scala 136:19]
  wire [3:0] _GEN_61 = _T_29 ? 4'h8 : _GEN_55; // @[Conditional.scala 39:67 ctrl.scala 137:20]
  wire [3:0] _GEN_62 = _T_29 ? 4'h5 : _GEN_56; // @[Conditional.scala 39:67 ctrl.scala 138:19]
  wire [2:0] _GEN_63 = _T_29 ? 3'h4 : {{1'd0}, _GEN_57}; // @[Conditional.scala 39:67 ctrl.scala 139:18]
  wire [3:0] _GEN_64 = _T_29 ? 4'h4 : _GEN_58; // @[Conditional.scala 39:67 ctrl.scala 140:19]
  wire [3:0] _GEN_65 = _T_22 ? 4'h0 : _GEN_60; // @[Conditional.scala 39:67 ctrl.scala 112:19]
  wire [3:0] _GEN_66 = _T_22 ? 4'h4 : _GEN_62; // @[Conditional.scala 39:67 ctrl.scala 113:19]
  wire [2:0] _GEN_67 = _T_22 ? 3'h0 : _GEN_63; // @[Conditional.scala 39:67 ctrl.scala 114:18]
  wire [3:0] _GEN_68 = _T_22 ? 4'h3 : _GEN_64; // @[Conditional.scala 39:67 ctrl.scala 115:19]
  wire [3:0] _GEN_69 = _T_22 ? {{1'd0}, _GEN_27} : _GEN_61; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_70 = _T_21 ? 4'h0 : _GEN_65; // @[Conditional.scala 39:67 ctrl.scala 104:19]
  wire [3:0] _GEN_71 = _T_21 ? 4'h2 : _GEN_69; // @[Conditional.scala 39:67 ctrl.scala 105:20]
  wire [3:0] _GEN_72 = _T_21 ? 4'h3 : _GEN_66; // @[Conditional.scala 39:67 ctrl.scala 106:19]
  wire [2:0] _GEN_73 = _T_21 ? 3'h2 : _GEN_67; // @[Conditional.scala 39:67 ctrl.scala 107:18]
  wire [3:0] _GEN_74 = _T_21 ? 4'h2 : _GEN_68; // @[Conditional.scala 39:67 ctrl.scala 108:19]
  wire [3:0] _GEN_75 = _T_9 ? 4'h0 : _GEN_71; // @[Conditional.scala 39:67 ctrl.scala 57:22]
  wire [2:0] _GEN_76 = _T_9 ? 3'h0 : _GEN_73; // @[Conditional.scala 39:67 ctrl.scala 58:22]
  wire [3:0] _GEN_77 = _T_9 ? 4'h0 : _GEN_74; // @[Conditional.scala 39:67 ctrl.scala 59:22]
  wire [3:0] _GEN_78 = _T_9 ? _GEN_21 : _GEN_70; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_79 = _T_9 ? {{2'd0}, _GEN_22} : _GEN_72; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_80 = _T_1 ? 4'h1 : _GEN_75; // @[Conditional.scala 40:58 ctrl.scala 29:22]
  wire [3:0] _GEN_81 = _T_1 ? 4'h1 : _GEN_79; // @[Conditional.scala 40:58 ctrl.scala 30:22]
  wire [2:0] _GEN_82 = _T_1 ? 3'h1 : _GEN_76; // @[Conditional.scala 40:58 ctrl.scala 31:22]
  wire [3:0] _GEN_83 = _T_1 ? 4'h1 : _GEN_77; // @[Conditional.scala 40:58 ctrl.scala 32:22]
  wire [3:0] _GEN_84 = _T_1 ? _GEN_5 : _GEN_78; // @[Conditional.scala 40:58]
  assign io_pc_ctrl = {{5'd0}, _GEN_82}; // @[Conditional.scala 40:58 ctrl.scala 31:22]
  assign io_imm_ctrl = {{4'd0}, _GEN_81}; // @[Conditional.scala 40:58 ctrl.scala 30:22]
  assign io_data_ctrl = {{4'd0}, _GEN_80}; // @[Conditional.scala 40:58 ctrl.scala 29:22]
  assign io_select_ctrl = {{4'd0}, _GEN_83}; // @[Conditional.scala 40:58 ctrl.scala 32:22]
  assign io_reg_ctrl = {{4'd0}, _GEN_83}; // @[Conditional.scala 40:58 ctrl.scala 32:22]
  assign io_alu_ctrl = {{4'd0}, _GEN_84}; // @[Conditional.scala 40:58]
endmodule
module data(
  input         clock,
  input         reset,
  input  [7:0]  io_data_ctrl,
  input  [31:0] io_data_addr,
  input  [31:0] io_data_write,
  output [31:0] io_data_read
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0; // @[data.scala 18:16]
  reg [31:0] mem_1; // @[data.scala 18:16]
  reg [31:0] mem_2; // @[data.scala 18:16]
  reg [31:0] mem_3; // @[data.scala 18:16]
  reg [31:0] mem_4; // @[data.scala 18:16]
  reg [31:0] mem_5; // @[data.scala 18:16]
  reg [31:0] mem_6; // @[data.scala 18:16]
  reg [31:0] mem_7; // @[data.scala 18:16]
  reg [31:0] mem_8; // @[data.scala 18:16]
  reg [31:0] mem_9; // @[data.scala 18:16]
  reg [31:0] mem_10; // @[data.scala 18:16]
  reg [31:0] mem_11; // @[data.scala 18:16]
  reg [31:0] mem_12; // @[data.scala 18:16]
  reg [31:0] mem_13; // @[data.scala 18:16]
  reg [31:0] mem_14; // @[data.scala 18:16]
  reg [31:0] mem_15; // @[data.scala 18:16]
  reg [31:0] mem_16; // @[data.scala 18:16]
  reg [31:0] mem_17; // @[data.scala 18:16]
  reg [31:0] mem_18; // @[data.scala 18:16]
  reg [31:0] mem_19; // @[data.scala 18:16]
  reg [31:0] mem_20; // @[data.scala 18:16]
  reg [31:0] mem_21; // @[data.scala 18:16]
  reg [31:0] mem_22; // @[data.scala 18:16]
  reg [31:0] mem_23; // @[data.scala 18:16]
  reg [31:0] mem_24; // @[data.scala 18:16]
  reg [31:0] mem_25; // @[data.scala 18:16]
  reg [31:0] mem_26; // @[data.scala 18:16]
  reg [31:0] mem_27; // @[data.scala 18:16]
  reg [31:0] mem_28; // @[data.scala 18:16]
  reg [31:0] mem_29; // @[data.scala 18:16]
  reg [31:0] mem_30; // @[data.scala 18:16]
  reg [31:0] mem_31; // @[data.scala 18:16]
  reg [31:0] mem_32; // @[data.scala 18:16]
  reg [31:0] mem_33; // @[data.scala 18:16]
  reg [31:0] mem_34; // @[data.scala 18:16]
  reg [31:0] mem_35; // @[data.scala 18:16]
  reg [31:0] mem_36; // @[data.scala 18:16]
  reg [31:0] mem_37; // @[data.scala 18:16]
  reg [31:0] mem_38; // @[data.scala 18:16]
  reg [31:0] mem_39; // @[data.scala 18:16]
  reg [31:0] mem_40; // @[data.scala 18:16]
  reg [31:0] mem_41; // @[data.scala 18:16]
  reg [31:0] mem_42; // @[data.scala 18:16]
  reg [31:0] mem_43; // @[data.scala 18:16]
  reg [31:0] mem_44; // @[data.scala 18:16]
  reg [31:0] mem_45; // @[data.scala 18:16]
  reg [31:0] mem_46; // @[data.scala 18:16]
  reg [31:0] mem_47; // @[data.scala 18:16]
  reg [31:0] mem_48; // @[data.scala 18:16]
  reg [31:0] mem_49; // @[data.scala 18:16]
  reg [31:0] mem_50; // @[data.scala 18:16]
  reg [31:0] mem_51; // @[data.scala 18:16]
  reg [31:0] mem_52; // @[data.scala 18:16]
  reg [31:0] mem_53; // @[data.scala 18:16]
  reg [31:0] mem_54; // @[data.scala 18:16]
  reg [31:0] mem_55; // @[data.scala 18:16]
  reg [31:0] mem_56; // @[data.scala 18:16]
  reg [31:0] mem_57; // @[data.scala 18:16]
  reg [31:0] mem_58; // @[data.scala 18:16]
  reg [31:0] mem_59; // @[data.scala 18:16]
  reg [31:0] mem_60; // @[data.scala 18:16]
  reg [31:0] mem_61; // @[data.scala 18:16]
  reg [31:0] mem_62; // @[data.scala 18:16]
  reg [31:0] mem_63; // @[data.scala 18:16]
  reg [31:0] mem_64; // @[data.scala 18:16]
  reg [31:0] mem_65; // @[data.scala 18:16]
  reg [31:0] mem_66; // @[data.scala 18:16]
  reg [31:0] mem_67; // @[data.scala 18:16]
  reg [31:0] mem_68; // @[data.scala 18:16]
  reg [31:0] mem_69; // @[data.scala 18:16]
  reg [31:0] mem_70; // @[data.scala 18:16]
  reg [31:0] mem_71; // @[data.scala 18:16]
  reg [31:0] mem_72; // @[data.scala 18:16]
  reg [31:0] mem_73; // @[data.scala 18:16]
  reg [31:0] mem_74; // @[data.scala 18:16]
  reg [31:0] mem_75; // @[data.scala 18:16]
  reg [31:0] mem_76; // @[data.scala 18:16]
  reg [31:0] mem_77; // @[data.scala 18:16]
  reg [31:0] mem_78; // @[data.scala 18:16]
  reg [31:0] mem_79; // @[data.scala 18:16]
  reg [31:0] mem_80; // @[data.scala 18:16]
  reg [31:0] mem_81; // @[data.scala 18:16]
  reg [31:0] mem_82; // @[data.scala 18:16]
  reg [31:0] mem_83; // @[data.scala 18:16]
  reg [31:0] mem_84; // @[data.scala 18:16]
  reg [31:0] mem_85; // @[data.scala 18:16]
  reg [31:0] mem_86; // @[data.scala 18:16]
  reg [31:0] mem_87; // @[data.scala 18:16]
  reg [31:0] mem_88; // @[data.scala 18:16]
  reg [31:0] mem_89; // @[data.scala 18:16]
  reg [31:0] mem_90; // @[data.scala 18:16]
  reg [31:0] mem_91; // @[data.scala 18:16]
  reg [31:0] mem_92; // @[data.scala 18:16]
  reg [31:0] mem_93; // @[data.scala 18:16]
  reg [31:0] mem_94; // @[data.scala 18:16]
  reg [31:0] mem_95; // @[data.scala 18:16]
  reg [31:0] mem_96; // @[data.scala 18:16]
  reg [31:0] mem_97; // @[data.scala 18:16]
  reg [31:0] mem_98; // @[data.scala 18:16]
  reg [31:0] mem_99; // @[data.scala 18:16]
  reg [31:0] mem_100; // @[data.scala 18:16]
  reg [31:0] mem_101; // @[data.scala 18:16]
  reg [31:0] mem_102; // @[data.scala 18:16]
  reg [31:0] mem_103; // @[data.scala 18:16]
  reg [31:0] mem_104; // @[data.scala 18:16]
  reg [31:0] mem_105; // @[data.scala 18:16]
  reg [31:0] mem_106; // @[data.scala 18:16]
  reg [31:0] mem_107; // @[data.scala 18:16]
  reg [31:0] mem_108; // @[data.scala 18:16]
  reg [31:0] mem_109; // @[data.scala 18:16]
  reg [31:0] mem_110; // @[data.scala 18:16]
  reg [31:0] mem_111; // @[data.scala 18:16]
  reg [31:0] mem_112; // @[data.scala 18:16]
  reg [31:0] mem_113; // @[data.scala 18:16]
  reg [31:0] mem_114; // @[data.scala 18:16]
  reg [31:0] mem_115; // @[data.scala 18:16]
  reg [31:0] mem_116; // @[data.scala 18:16]
  reg [31:0] mem_117; // @[data.scala 18:16]
  reg [31:0] mem_118; // @[data.scala 18:16]
  reg [31:0] mem_119; // @[data.scala 18:16]
  reg [31:0] mem_120; // @[data.scala 18:16]
  reg [31:0] mem_121; // @[data.scala 18:16]
  reg [31:0] mem_122; // @[data.scala 18:16]
  reg [31:0] mem_123; // @[data.scala 18:16]
  reg [31:0] mem_124; // @[data.scala 18:16]
  reg [31:0] mem_125; // @[data.scala 18:16]
  reg [31:0] mem_126; // @[data.scala 18:16]
  reg [31:0] mem_127; // @[data.scala 18:16]
  wire  _T_1 = 8'hd == io_data_ctrl; // @[Conditional.scala 37:30]
  wire  _T_2 = 8'h1 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire  _T_3 = 8'h0 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire  _T_4 = 8'h8 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire  _T_5 = 8'h2 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire  _T_6 = 8'h3 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_1 = 7'h1 == io_data_addr[6:0] ? mem_1 : mem_0; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_2 = 7'h2 == io_data_addr[6:0] ? mem_2 : _GEN_1; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_3 = 7'h3 == io_data_addr[6:0] ? mem_3 : _GEN_2; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_4 = 7'h4 == io_data_addr[6:0] ? mem_4 : _GEN_3; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_5 = 7'h5 == io_data_addr[6:0] ? mem_5 : _GEN_4; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_6 = 7'h6 == io_data_addr[6:0] ? mem_6 : _GEN_5; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_7 = 7'h7 == io_data_addr[6:0] ? mem_7 : _GEN_6; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_8 = 7'h8 == io_data_addr[6:0] ? mem_8 : _GEN_7; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_9 = 7'h9 == io_data_addr[6:0] ? mem_9 : _GEN_8; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_10 = 7'ha == io_data_addr[6:0] ? mem_10 : _GEN_9; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_11 = 7'hb == io_data_addr[6:0] ? mem_11 : _GEN_10; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_12 = 7'hc == io_data_addr[6:0] ? mem_12 : _GEN_11; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_13 = 7'hd == io_data_addr[6:0] ? mem_13 : _GEN_12; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_14 = 7'he == io_data_addr[6:0] ? mem_14 : _GEN_13; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_15 = 7'hf == io_data_addr[6:0] ? mem_15 : _GEN_14; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_16 = 7'h10 == io_data_addr[6:0] ? mem_16 : _GEN_15; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_17 = 7'h11 == io_data_addr[6:0] ? mem_17 : _GEN_16; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_18 = 7'h12 == io_data_addr[6:0] ? mem_18 : _GEN_17; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_19 = 7'h13 == io_data_addr[6:0] ? mem_19 : _GEN_18; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_20 = 7'h14 == io_data_addr[6:0] ? mem_20 : _GEN_19; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_21 = 7'h15 == io_data_addr[6:0] ? mem_21 : _GEN_20; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_22 = 7'h16 == io_data_addr[6:0] ? mem_22 : _GEN_21; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_23 = 7'h17 == io_data_addr[6:0] ? mem_23 : _GEN_22; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_24 = 7'h18 == io_data_addr[6:0] ? mem_24 : _GEN_23; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_25 = 7'h19 == io_data_addr[6:0] ? mem_25 : _GEN_24; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_26 = 7'h1a == io_data_addr[6:0] ? mem_26 : _GEN_25; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_27 = 7'h1b == io_data_addr[6:0] ? mem_27 : _GEN_26; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_28 = 7'h1c == io_data_addr[6:0] ? mem_28 : _GEN_27; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_29 = 7'h1d == io_data_addr[6:0] ? mem_29 : _GEN_28; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_30 = 7'h1e == io_data_addr[6:0] ? mem_30 : _GEN_29; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_31 = 7'h1f == io_data_addr[6:0] ? mem_31 : _GEN_30; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_32 = 7'h20 == io_data_addr[6:0] ? mem_32 : _GEN_31; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_33 = 7'h21 == io_data_addr[6:0] ? mem_33 : _GEN_32; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_34 = 7'h22 == io_data_addr[6:0] ? mem_34 : _GEN_33; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_35 = 7'h23 == io_data_addr[6:0] ? mem_35 : _GEN_34; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_36 = 7'h24 == io_data_addr[6:0] ? mem_36 : _GEN_35; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_37 = 7'h25 == io_data_addr[6:0] ? mem_37 : _GEN_36; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_38 = 7'h26 == io_data_addr[6:0] ? mem_38 : _GEN_37; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_39 = 7'h27 == io_data_addr[6:0] ? mem_39 : _GEN_38; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_40 = 7'h28 == io_data_addr[6:0] ? mem_40 : _GEN_39; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_41 = 7'h29 == io_data_addr[6:0] ? mem_41 : _GEN_40; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_42 = 7'h2a == io_data_addr[6:0] ? mem_42 : _GEN_41; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_43 = 7'h2b == io_data_addr[6:0] ? mem_43 : _GEN_42; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_44 = 7'h2c == io_data_addr[6:0] ? mem_44 : _GEN_43; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_45 = 7'h2d == io_data_addr[6:0] ? mem_45 : _GEN_44; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_46 = 7'h2e == io_data_addr[6:0] ? mem_46 : _GEN_45; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_47 = 7'h2f == io_data_addr[6:0] ? mem_47 : _GEN_46; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_48 = 7'h30 == io_data_addr[6:0] ? mem_48 : _GEN_47; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_49 = 7'h31 == io_data_addr[6:0] ? mem_49 : _GEN_48; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_50 = 7'h32 == io_data_addr[6:0] ? mem_50 : _GEN_49; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_51 = 7'h33 == io_data_addr[6:0] ? mem_51 : _GEN_50; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_52 = 7'h34 == io_data_addr[6:0] ? mem_52 : _GEN_51; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_53 = 7'h35 == io_data_addr[6:0] ? mem_53 : _GEN_52; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_54 = 7'h36 == io_data_addr[6:0] ? mem_54 : _GEN_53; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_55 = 7'h37 == io_data_addr[6:0] ? mem_55 : _GEN_54; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_56 = 7'h38 == io_data_addr[6:0] ? mem_56 : _GEN_55; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_57 = 7'h39 == io_data_addr[6:0] ? mem_57 : _GEN_56; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_58 = 7'h3a == io_data_addr[6:0] ? mem_58 : _GEN_57; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_59 = 7'h3b == io_data_addr[6:0] ? mem_59 : _GEN_58; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_60 = 7'h3c == io_data_addr[6:0] ? mem_60 : _GEN_59; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_61 = 7'h3d == io_data_addr[6:0] ? mem_61 : _GEN_60; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_62 = 7'h3e == io_data_addr[6:0] ? mem_62 : _GEN_61; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_63 = 7'h3f == io_data_addr[6:0] ? mem_63 : _GEN_62; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_64 = 7'h40 == io_data_addr[6:0] ? mem_64 : _GEN_63; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_65 = 7'h41 == io_data_addr[6:0] ? mem_65 : _GEN_64; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_66 = 7'h42 == io_data_addr[6:0] ? mem_66 : _GEN_65; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_67 = 7'h43 == io_data_addr[6:0] ? mem_67 : _GEN_66; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_68 = 7'h44 == io_data_addr[6:0] ? mem_68 : _GEN_67; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_69 = 7'h45 == io_data_addr[6:0] ? mem_69 : _GEN_68; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_70 = 7'h46 == io_data_addr[6:0] ? mem_70 : _GEN_69; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_71 = 7'h47 == io_data_addr[6:0] ? mem_71 : _GEN_70; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_72 = 7'h48 == io_data_addr[6:0] ? mem_72 : _GEN_71; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_73 = 7'h49 == io_data_addr[6:0] ? mem_73 : _GEN_72; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_74 = 7'h4a == io_data_addr[6:0] ? mem_74 : _GEN_73; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_75 = 7'h4b == io_data_addr[6:0] ? mem_75 : _GEN_74; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_76 = 7'h4c == io_data_addr[6:0] ? mem_76 : _GEN_75; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_77 = 7'h4d == io_data_addr[6:0] ? mem_77 : _GEN_76; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_78 = 7'h4e == io_data_addr[6:0] ? mem_78 : _GEN_77; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_79 = 7'h4f == io_data_addr[6:0] ? mem_79 : _GEN_78; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_80 = 7'h50 == io_data_addr[6:0] ? mem_80 : _GEN_79; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_81 = 7'h51 == io_data_addr[6:0] ? mem_81 : _GEN_80; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_82 = 7'h52 == io_data_addr[6:0] ? mem_82 : _GEN_81; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_83 = 7'h53 == io_data_addr[6:0] ? mem_83 : _GEN_82; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_84 = 7'h54 == io_data_addr[6:0] ? mem_84 : _GEN_83; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_85 = 7'h55 == io_data_addr[6:0] ? mem_85 : _GEN_84; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_86 = 7'h56 == io_data_addr[6:0] ? mem_86 : _GEN_85; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_87 = 7'h57 == io_data_addr[6:0] ? mem_87 : _GEN_86; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_88 = 7'h58 == io_data_addr[6:0] ? mem_88 : _GEN_87; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_89 = 7'h59 == io_data_addr[6:0] ? mem_89 : _GEN_88; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_90 = 7'h5a == io_data_addr[6:0] ? mem_90 : _GEN_89; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_91 = 7'h5b == io_data_addr[6:0] ? mem_91 : _GEN_90; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_92 = 7'h5c == io_data_addr[6:0] ? mem_92 : _GEN_91; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_93 = 7'h5d == io_data_addr[6:0] ? mem_93 : _GEN_92; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_94 = 7'h5e == io_data_addr[6:0] ? mem_94 : _GEN_93; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_95 = 7'h5f == io_data_addr[6:0] ? mem_95 : _GEN_94; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_96 = 7'h60 == io_data_addr[6:0] ? mem_96 : _GEN_95; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_97 = 7'h61 == io_data_addr[6:0] ? mem_97 : _GEN_96; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_98 = 7'h62 == io_data_addr[6:0] ? mem_98 : _GEN_97; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_99 = 7'h63 == io_data_addr[6:0] ? mem_99 : _GEN_98; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_100 = 7'h64 == io_data_addr[6:0] ? mem_100 : _GEN_99; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_101 = 7'h65 == io_data_addr[6:0] ? mem_101 : _GEN_100; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_102 = 7'h66 == io_data_addr[6:0] ? mem_102 : _GEN_101; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_103 = 7'h67 == io_data_addr[6:0] ? mem_103 : _GEN_102; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_104 = 7'h68 == io_data_addr[6:0] ? mem_104 : _GEN_103; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_105 = 7'h69 == io_data_addr[6:0] ? mem_105 : _GEN_104; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_106 = 7'h6a == io_data_addr[6:0] ? mem_106 : _GEN_105; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_107 = 7'h6b == io_data_addr[6:0] ? mem_107 : _GEN_106; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_108 = 7'h6c == io_data_addr[6:0] ? mem_108 : _GEN_107; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_109 = 7'h6d == io_data_addr[6:0] ? mem_109 : _GEN_108; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_110 = 7'h6e == io_data_addr[6:0] ? mem_110 : _GEN_109; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_111 = 7'h6f == io_data_addr[6:0] ? mem_111 : _GEN_110; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_112 = 7'h70 == io_data_addr[6:0] ? mem_112 : _GEN_111; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_113 = 7'h71 == io_data_addr[6:0] ? mem_113 : _GEN_112; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_114 = 7'h72 == io_data_addr[6:0] ? mem_114 : _GEN_113; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_115 = 7'h73 == io_data_addr[6:0] ? mem_115 : _GEN_114; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_116 = 7'h74 == io_data_addr[6:0] ? mem_116 : _GEN_115; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_117 = 7'h75 == io_data_addr[6:0] ? mem_117 : _GEN_116; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_118 = 7'h76 == io_data_addr[6:0] ? mem_118 : _GEN_117; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_119 = 7'h77 == io_data_addr[6:0] ? mem_119 : _GEN_118; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_120 = 7'h78 == io_data_addr[6:0] ? mem_120 : _GEN_119; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_121 = 7'h79 == io_data_addr[6:0] ? mem_121 : _GEN_120; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_122 = 7'h7a == io_data_addr[6:0] ? mem_122 : _GEN_121; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_123 = 7'h7b == io_data_addr[6:0] ? mem_123 : _GEN_122; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_124 = 7'h7c == io_data_addr[6:0] ? mem_124 : _GEN_123; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_125 = 7'h7d == io_data_addr[6:0] ? mem_125 : _GEN_124; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_126 = 7'h7e == io_data_addr[6:0] ? mem_126 : _GEN_125; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_127 = 7'h7f == io_data_addr[6:0] ? mem_127 : _GEN_126; // @[data.scala 44:29 data.scala 44:29]
  wire [31:0] _GEN_3730 = {{24'd0}, _GEN_127[7:0]}; // @[data.scala 45:48]
  wire [31:0] _io_data_read_T_3 = _GEN_3730 + 32'hffffff00; // @[data.scala 45:48]
  wire [31:0] _GEN_384 = _GEN_127[7] ? _io_data_read_T_3 : {{24'd0}, _GEN_127[7:0]}; // @[data.scala 44:41 data.scala 45:22 data.scala 48:22]
  wire  _T_10 = 8'h6 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire  _T_11 = 8'h4 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_3731 = {{16'd0}, _GEN_127[15:0]}; // @[data.scala 56:49]
  wire [31:0] _io_data_read_T_11 = _GEN_3731 + 32'hffff0000; // @[data.scala 56:49]
  wire [31:0] _GEN_897 = _GEN_127[15] ? _io_data_read_T_11 : {{16'd0}, _GEN_127[15:0]}; // @[data.scala 55:42 data.scala 56:22 data.scala 59:22]
  wire  _T_15 = 8'h7 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire  _T_16 = 8'he == io_data_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _io_data_read_T_18 = {_GEN_127[31:12], 12'h0}; // @[data.scala 66:48]
  wire  _T_17 = 8'h5 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire  _T_18 = 8'h9 == io_data_ctrl; // @[Conditional.scala 37:30]
  wire  _T_19 = 8'ha == io_data_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _mem_T_20 = {{24'd0}, io_data_write[7:0]}; // @[data.scala 76:25 data.scala 76:25]
  wire [31:0] _GEN_1282 = 7'h0 == io_data_addr[6:0] ? _mem_T_20 : mem_0; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1283 = 7'h1 == io_data_addr[6:0] ? _mem_T_20 : mem_1; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1284 = 7'h2 == io_data_addr[6:0] ? _mem_T_20 : mem_2; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1285 = 7'h3 == io_data_addr[6:0] ? _mem_T_20 : mem_3; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1286 = 7'h4 == io_data_addr[6:0] ? _mem_T_20 : mem_4; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1287 = 7'h5 == io_data_addr[6:0] ? _mem_T_20 : mem_5; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1288 = 7'h6 == io_data_addr[6:0] ? _mem_T_20 : mem_6; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1289 = 7'h7 == io_data_addr[6:0] ? _mem_T_20 : mem_7; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1290 = 7'h8 == io_data_addr[6:0] ? _mem_T_20 : mem_8; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1291 = 7'h9 == io_data_addr[6:0] ? _mem_T_20 : mem_9; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1292 = 7'ha == io_data_addr[6:0] ? _mem_T_20 : mem_10; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1293 = 7'hb == io_data_addr[6:0] ? _mem_T_20 : mem_11; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1294 = 7'hc == io_data_addr[6:0] ? _mem_T_20 : mem_12; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1295 = 7'hd == io_data_addr[6:0] ? _mem_T_20 : mem_13; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1296 = 7'he == io_data_addr[6:0] ? _mem_T_20 : mem_14; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1297 = 7'hf == io_data_addr[6:0] ? _mem_T_20 : mem_15; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1298 = 7'h10 == io_data_addr[6:0] ? _mem_T_20 : mem_16; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1299 = 7'h11 == io_data_addr[6:0] ? _mem_T_20 : mem_17; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1300 = 7'h12 == io_data_addr[6:0] ? _mem_T_20 : mem_18; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1301 = 7'h13 == io_data_addr[6:0] ? _mem_T_20 : mem_19; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1302 = 7'h14 == io_data_addr[6:0] ? _mem_T_20 : mem_20; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1303 = 7'h15 == io_data_addr[6:0] ? _mem_T_20 : mem_21; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1304 = 7'h16 == io_data_addr[6:0] ? _mem_T_20 : mem_22; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1305 = 7'h17 == io_data_addr[6:0] ? _mem_T_20 : mem_23; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1306 = 7'h18 == io_data_addr[6:0] ? _mem_T_20 : mem_24; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1307 = 7'h19 == io_data_addr[6:0] ? _mem_T_20 : mem_25; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1308 = 7'h1a == io_data_addr[6:0] ? _mem_T_20 : mem_26; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1309 = 7'h1b == io_data_addr[6:0] ? _mem_T_20 : mem_27; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1310 = 7'h1c == io_data_addr[6:0] ? _mem_T_20 : mem_28; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1311 = 7'h1d == io_data_addr[6:0] ? _mem_T_20 : mem_29; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1312 = 7'h1e == io_data_addr[6:0] ? _mem_T_20 : mem_30; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1313 = 7'h1f == io_data_addr[6:0] ? _mem_T_20 : mem_31; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1314 = 7'h20 == io_data_addr[6:0] ? _mem_T_20 : mem_32; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1315 = 7'h21 == io_data_addr[6:0] ? _mem_T_20 : mem_33; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1316 = 7'h22 == io_data_addr[6:0] ? _mem_T_20 : mem_34; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1317 = 7'h23 == io_data_addr[6:0] ? _mem_T_20 : mem_35; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1318 = 7'h24 == io_data_addr[6:0] ? _mem_T_20 : mem_36; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1319 = 7'h25 == io_data_addr[6:0] ? _mem_T_20 : mem_37; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1320 = 7'h26 == io_data_addr[6:0] ? _mem_T_20 : mem_38; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1321 = 7'h27 == io_data_addr[6:0] ? _mem_T_20 : mem_39; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1322 = 7'h28 == io_data_addr[6:0] ? _mem_T_20 : mem_40; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1323 = 7'h29 == io_data_addr[6:0] ? _mem_T_20 : mem_41; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1324 = 7'h2a == io_data_addr[6:0] ? _mem_T_20 : mem_42; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1325 = 7'h2b == io_data_addr[6:0] ? _mem_T_20 : mem_43; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1326 = 7'h2c == io_data_addr[6:0] ? _mem_T_20 : mem_44; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1327 = 7'h2d == io_data_addr[6:0] ? _mem_T_20 : mem_45; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1328 = 7'h2e == io_data_addr[6:0] ? _mem_T_20 : mem_46; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1329 = 7'h2f == io_data_addr[6:0] ? _mem_T_20 : mem_47; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1330 = 7'h30 == io_data_addr[6:0] ? _mem_T_20 : mem_48; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1331 = 7'h31 == io_data_addr[6:0] ? _mem_T_20 : mem_49; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1332 = 7'h32 == io_data_addr[6:0] ? _mem_T_20 : mem_50; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1333 = 7'h33 == io_data_addr[6:0] ? _mem_T_20 : mem_51; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1334 = 7'h34 == io_data_addr[6:0] ? _mem_T_20 : mem_52; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1335 = 7'h35 == io_data_addr[6:0] ? _mem_T_20 : mem_53; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1336 = 7'h36 == io_data_addr[6:0] ? _mem_T_20 : mem_54; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1337 = 7'h37 == io_data_addr[6:0] ? _mem_T_20 : mem_55; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1338 = 7'h38 == io_data_addr[6:0] ? _mem_T_20 : mem_56; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1339 = 7'h39 == io_data_addr[6:0] ? _mem_T_20 : mem_57; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1340 = 7'h3a == io_data_addr[6:0] ? _mem_T_20 : mem_58; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1341 = 7'h3b == io_data_addr[6:0] ? _mem_T_20 : mem_59; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1342 = 7'h3c == io_data_addr[6:0] ? _mem_T_20 : mem_60; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1343 = 7'h3d == io_data_addr[6:0] ? _mem_T_20 : mem_61; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1344 = 7'h3e == io_data_addr[6:0] ? _mem_T_20 : mem_62; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1345 = 7'h3f == io_data_addr[6:0] ? _mem_T_20 : mem_63; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1346 = 7'h40 == io_data_addr[6:0] ? _mem_T_20 : mem_64; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1347 = 7'h41 == io_data_addr[6:0] ? _mem_T_20 : mem_65; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1348 = 7'h42 == io_data_addr[6:0] ? _mem_T_20 : mem_66; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1349 = 7'h43 == io_data_addr[6:0] ? _mem_T_20 : mem_67; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1350 = 7'h44 == io_data_addr[6:0] ? _mem_T_20 : mem_68; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1351 = 7'h45 == io_data_addr[6:0] ? _mem_T_20 : mem_69; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1352 = 7'h46 == io_data_addr[6:0] ? _mem_T_20 : mem_70; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1353 = 7'h47 == io_data_addr[6:0] ? _mem_T_20 : mem_71; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1354 = 7'h48 == io_data_addr[6:0] ? _mem_T_20 : mem_72; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1355 = 7'h49 == io_data_addr[6:0] ? _mem_T_20 : mem_73; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1356 = 7'h4a == io_data_addr[6:0] ? _mem_T_20 : mem_74; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1357 = 7'h4b == io_data_addr[6:0] ? _mem_T_20 : mem_75; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1358 = 7'h4c == io_data_addr[6:0] ? _mem_T_20 : mem_76; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1359 = 7'h4d == io_data_addr[6:0] ? _mem_T_20 : mem_77; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1360 = 7'h4e == io_data_addr[6:0] ? _mem_T_20 : mem_78; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1361 = 7'h4f == io_data_addr[6:0] ? _mem_T_20 : mem_79; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1362 = 7'h50 == io_data_addr[6:0] ? _mem_T_20 : mem_80; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1363 = 7'h51 == io_data_addr[6:0] ? _mem_T_20 : mem_81; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1364 = 7'h52 == io_data_addr[6:0] ? _mem_T_20 : mem_82; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1365 = 7'h53 == io_data_addr[6:0] ? _mem_T_20 : mem_83; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1366 = 7'h54 == io_data_addr[6:0] ? _mem_T_20 : mem_84; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1367 = 7'h55 == io_data_addr[6:0] ? _mem_T_20 : mem_85; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1368 = 7'h56 == io_data_addr[6:0] ? _mem_T_20 : mem_86; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1369 = 7'h57 == io_data_addr[6:0] ? _mem_T_20 : mem_87; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1370 = 7'h58 == io_data_addr[6:0] ? _mem_T_20 : mem_88; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1371 = 7'h59 == io_data_addr[6:0] ? _mem_T_20 : mem_89; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1372 = 7'h5a == io_data_addr[6:0] ? _mem_T_20 : mem_90; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1373 = 7'h5b == io_data_addr[6:0] ? _mem_T_20 : mem_91; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1374 = 7'h5c == io_data_addr[6:0] ? _mem_T_20 : mem_92; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1375 = 7'h5d == io_data_addr[6:0] ? _mem_T_20 : mem_93; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1376 = 7'h5e == io_data_addr[6:0] ? _mem_T_20 : mem_94; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1377 = 7'h5f == io_data_addr[6:0] ? _mem_T_20 : mem_95; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1378 = 7'h60 == io_data_addr[6:0] ? _mem_T_20 : mem_96; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1379 = 7'h61 == io_data_addr[6:0] ? _mem_T_20 : mem_97; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1380 = 7'h62 == io_data_addr[6:0] ? _mem_T_20 : mem_98; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1381 = 7'h63 == io_data_addr[6:0] ? _mem_T_20 : mem_99; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1382 = 7'h64 == io_data_addr[6:0] ? _mem_T_20 : mem_100; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1383 = 7'h65 == io_data_addr[6:0] ? _mem_T_20 : mem_101; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1384 = 7'h66 == io_data_addr[6:0] ? _mem_T_20 : mem_102; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1385 = 7'h67 == io_data_addr[6:0] ? _mem_T_20 : mem_103; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1386 = 7'h68 == io_data_addr[6:0] ? _mem_T_20 : mem_104; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1387 = 7'h69 == io_data_addr[6:0] ? _mem_T_20 : mem_105; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1388 = 7'h6a == io_data_addr[6:0] ? _mem_T_20 : mem_106; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1389 = 7'h6b == io_data_addr[6:0] ? _mem_T_20 : mem_107; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1390 = 7'h6c == io_data_addr[6:0] ? _mem_T_20 : mem_108; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1391 = 7'h6d == io_data_addr[6:0] ? _mem_T_20 : mem_109; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1392 = 7'h6e == io_data_addr[6:0] ? _mem_T_20 : mem_110; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1393 = 7'h6f == io_data_addr[6:0] ? _mem_T_20 : mem_111; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1394 = 7'h70 == io_data_addr[6:0] ? _mem_T_20 : mem_112; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1395 = 7'h71 == io_data_addr[6:0] ? _mem_T_20 : mem_113; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1396 = 7'h72 == io_data_addr[6:0] ? _mem_T_20 : mem_114; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1397 = 7'h73 == io_data_addr[6:0] ? _mem_T_20 : mem_115; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1398 = 7'h74 == io_data_addr[6:0] ? _mem_T_20 : mem_116; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1399 = 7'h75 == io_data_addr[6:0] ? _mem_T_20 : mem_117; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1400 = 7'h76 == io_data_addr[6:0] ? _mem_T_20 : mem_118; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1401 = 7'h77 == io_data_addr[6:0] ? _mem_T_20 : mem_119; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1402 = 7'h78 == io_data_addr[6:0] ? _mem_T_20 : mem_120; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1403 = 7'h79 == io_data_addr[6:0] ? _mem_T_20 : mem_121; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1404 = 7'h7a == io_data_addr[6:0] ? _mem_T_20 : mem_122; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1405 = 7'h7b == io_data_addr[6:0] ? _mem_T_20 : mem_123; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1406 = 7'h7c == io_data_addr[6:0] ? _mem_T_20 : mem_124; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1407 = 7'h7d == io_data_addr[6:0] ? _mem_T_20 : mem_125; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1408 = 7'h7e == io_data_addr[6:0] ? _mem_T_20 : mem_126; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire [31:0] _GEN_1409 = 7'h7f == io_data_addr[6:0] ? _mem_T_20 : mem_127; // @[data.scala 76:25 data.scala 76:25 data.scala 18:16]
  wire  _T_21 = 8'hb == io_data_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _mem_T_22 = {{16'd0}, io_data_write[15:0]}; // @[data.scala 80:25 data.scala 80:25]
  wire [31:0] _GEN_1410 = 7'h0 == io_data_addr[6:0] ? _mem_T_22 : mem_0; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1411 = 7'h1 == io_data_addr[6:0] ? _mem_T_22 : mem_1; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1412 = 7'h2 == io_data_addr[6:0] ? _mem_T_22 : mem_2; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1413 = 7'h3 == io_data_addr[6:0] ? _mem_T_22 : mem_3; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1414 = 7'h4 == io_data_addr[6:0] ? _mem_T_22 : mem_4; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1415 = 7'h5 == io_data_addr[6:0] ? _mem_T_22 : mem_5; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1416 = 7'h6 == io_data_addr[6:0] ? _mem_T_22 : mem_6; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1417 = 7'h7 == io_data_addr[6:0] ? _mem_T_22 : mem_7; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1418 = 7'h8 == io_data_addr[6:0] ? _mem_T_22 : mem_8; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1419 = 7'h9 == io_data_addr[6:0] ? _mem_T_22 : mem_9; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1420 = 7'ha == io_data_addr[6:0] ? _mem_T_22 : mem_10; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1421 = 7'hb == io_data_addr[6:0] ? _mem_T_22 : mem_11; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1422 = 7'hc == io_data_addr[6:0] ? _mem_T_22 : mem_12; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1423 = 7'hd == io_data_addr[6:0] ? _mem_T_22 : mem_13; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1424 = 7'he == io_data_addr[6:0] ? _mem_T_22 : mem_14; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1425 = 7'hf == io_data_addr[6:0] ? _mem_T_22 : mem_15; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1426 = 7'h10 == io_data_addr[6:0] ? _mem_T_22 : mem_16; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1427 = 7'h11 == io_data_addr[6:0] ? _mem_T_22 : mem_17; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1428 = 7'h12 == io_data_addr[6:0] ? _mem_T_22 : mem_18; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1429 = 7'h13 == io_data_addr[6:0] ? _mem_T_22 : mem_19; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1430 = 7'h14 == io_data_addr[6:0] ? _mem_T_22 : mem_20; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1431 = 7'h15 == io_data_addr[6:0] ? _mem_T_22 : mem_21; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1432 = 7'h16 == io_data_addr[6:0] ? _mem_T_22 : mem_22; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1433 = 7'h17 == io_data_addr[6:0] ? _mem_T_22 : mem_23; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1434 = 7'h18 == io_data_addr[6:0] ? _mem_T_22 : mem_24; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1435 = 7'h19 == io_data_addr[6:0] ? _mem_T_22 : mem_25; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1436 = 7'h1a == io_data_addr[6:0] ? _mem_T_22 : mem_26; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1437 = 7'h1b == io_data_addr[6:0] ? _mem_T_22 : mem_27; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1438 = 7'h1c == io_data_addr[6:0] ? _mem_T_22 : mem_28; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1439 = 7'h1d == io_data_addr[6:0] ? _mem_T_22 : mem_29; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1440 = 7'h1e == io_data_addr[6:0] ? _mem_T_22 : mem_30; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1441 = 7'h1f == io_data_addr[6:0] ? _mem_T_22 : mem_31; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1442 = 7'h20 == io_data_addr[6:0] ? _mem_T_22 : mem_32; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1443 = 7'h21 == io_data_addr[6:0] ? _mem_T_22 : mem_33; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1444 = 7'h22 == io_data_addr[6:0] ? _mem_T_22 : mem_34; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1445 = 7'h23 == io_data_addr[6:0] ? _mem_T_22 : mem_35; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1446 = 7'h24 == io_data_addr[6:0] ? _mem_T_22 : mem_36; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1447 = 7'h25 == io_data_addr[6:0] ? _mem_T_22 : mem_37; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1448 = 7'h26 == io_data_addr[6:0] ? _mem_T_22 : mem_38; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1449 = 7'h27 == io_data_addr[6:0] ? _mem_T_22 : mem_39; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1450 = 7'h28 == io_data_addr[6:0] ? _mem_T_22 : mem_40; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1451 = 7'h29 == io_data_addr[6:0] ? _mem_T_22 : mem_41; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1452 = 7'h2a == io_data_addr[6:0] ? _mem_T_22 : mem_42; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1453 = 7'h2b == io_data_addr[6:0] ? _mem_T_22 : mem_43; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1454 = 7'h2c == io_data_addr[6:0] ? _mem_T_22 : mem_44; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1455 = 7'h2d == io_data_addr[6:0] ? _mem_T_22 : mem_45; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1456 = 7'h2e == io_data_addr[6:0] ? _mem_T_22 : mem_46; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1457 = 7'h2f == io_data_addr[6:0] ? _mem_T_22 : mem_47; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1458 = 7'h30 == io_data_addr[6:0] ? _mem_T_22 : mem_48; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1459 = 7'h31 == io_data_addr[6:0] ? _mem_T_22 : mem_49; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1460 = 7'h32 == io_data_addr[6:0] ? _mem_T_22 : mem_50; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1461 = 7'h33 == io_data_addr[6:0] ? _mem_T_22 : mem_51; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1462 = 7'h34 == io_data_addr[6:0] ? _mem_T_22 : mem_52; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1463 = 7'h35 == io_data_addr[6:0] ? _mem_T_22 : mem_53; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1464 = 7'h36 == io_data_addr[6:0] ? _mem_T_22 : mem_54; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1465 = 7'h37 == io_data_addr[6:0] ? _mem_T_22 : mem_55; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1466 = 7'h38 == io_data_addr[6:0] ? _mem_T_22 : mem_56; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1467 = 7'h39 == io_data_addr[6:0] ? _mem_T_22 : mem_57; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1468 = 7'h3a == io_data_addr[6:0] ? _mem_T_22 : mem_58; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1469 = 7'h3b == io_data_addr[6:0] ? _mem_T_22 : mem_59; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1470 = 7'h3c == io_data_addr[6:0] ? _mem_T_22 : mem_60; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1471 = 7'h3d == io_data_addr[6:0] ? _mem_T_22 : mem_61; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1472 = 7'h3e == io_data_addr[6:0] ? _mem_T_22 : mem_62; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1473 = 7'h3f == io_data_addr[6:0] ? _mem_T_22 : mem_63; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1474 = 7'h40 == io_data_addr[6:0] ? _mem_T_22 : mem_64; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1475 = 7'h41 == io_data_addr[6:0] ? _mem_T_22 : mem_65; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1476 = 7'h42 == io_data_addr[6:0] ? _mem_T_22 : mem_66; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1477 = 7'h43 == io_data_addr[6:0] ? _mem_T_22 : mem_67; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1478 = 7'h44 == io_data_addr[6:0] ? _mem_T_22 : mem_68; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1479 = 7'h45 == io_data_addr[6:0] ? _mem_T_22 : mem_69; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1480 = 7'h46 == io_data_addr[6:0] ? _mem_T_22 : mem_70; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1481 = 7'h47 == io_data_addr[6:0] ? _mem_T_22 : mem_71; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1482 = 7'h48 == io_data_addr[6:0] ? _mem_T_22 : mem_72; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1483 = 7'h49 == io_data_addr[6:0] ? _mem_T_22 : mem_73; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1484 = 7'h4a == io_data_addr[6:0] ? _mem_T_22 : mem_74; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1485 = 7'h4b == io_data_addr[6:0] ? _mem_T_22 : mem_75; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1486 = 7'h4c == io_data_addr[6:0] ? _mem_T_22 : mem_76; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1487 = 7'h4d == io_data_addr[6:0] ? _mem_T_22 : mem_77; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1488 = 7'h4e == io_data_addr[6:0] ? _mem_T_22 : mem_78; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1489 = 7'h4f == io_data_addr[6:0] ? _mem_T_22 : mem_79; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1490 = 7'h50 == io_data_addr[6:0] ? _mem_T_22 : mem_80; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1491 = 7'h51 == io_data_addr[6:0] ? _mem_T_22 : mem_81; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1492 = 7'h52 == io_data_addr[6:0] ? _mem_T_22 : mem_82; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1493 = 7'h53 == io_data_addr[6:0] ? _mem_T_22 : mem_83; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1494 = 7'h54 == io_data_addr[6:0] ? _mem_T_22 : mem_84; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1495 = 7'h55 == io_data_addr[6:0] ? _mem_T_22 : mem_85; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1496 = 7'h56 == io_data_addr[6:0] ? _mem_T_22 : mem_86; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1497 = 7'h57 == io_data_addr[6:0] ? _mem_T_22 : mem_87; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1498 = 7'h58 == io_data_addr[6:0] ? _mem_T_22 : mem_88; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1499 = 7'h59 == io_data_addr[6:0] ? _mem_T_22 : mem_89; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1500 = 7'h5a == io_data_addr[6:0] ? _mem_T_22 : mem_90; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1501 = 7'h5b == io_data_addr[6:0] ? _mem_T_22 : mem_91; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1502 = 7'h5c == io_data_addr[6:0] ? _mem_T_22 : mem_92; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1503 = 7'h5d == io_data_addr[6:0] ? _mem_T_22 : mem_93; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1504 = 7'h5e == io_data_addr[6:0] ? _mem_T_22 : mem_94; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1505 = 7'h5f == io_data_addr[6:0] ? _mem_T_22 : mem_95; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1506 = 7'h60 == io_data_addr[6:0] ? _mem_T_22 : mem_96; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1507 = 7'h61 == io_data_addr[6:0] ? _mem_T_22 : mem_97; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1508 = 7'h62 == io_data_addr[6:0] ? _mem_T_22 : mem_98; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1509 = 7'h63 == io_data_addr[6:0] ? _mem_T_22 : mem_99; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1510 = 7'h64 == io_data_addr[6:0] ? _mem_T_22 : mem_100; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1511 = 7'h65 == io_data_addr[6:0] ? _mem_T_22 : mem_101; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1512 = 7'h66 == io_data_addr[6:0] ? _mem_T_22 : mem_102; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1513 = 7'h67 == io_data_addr[6:0] ? _mem_T_22 : mem_103; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1514 = 7'h68 == io_data_addr[6:0] ? _mem_T_22 : mem_104; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1515 = 7'h69 == io_data_addr[6:0] ? _mem_T_22 : mem_105; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1516 = 7'h6a == io_data_addr[6:0] ? _mem_T_22 : mem_106; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1517 = 7'h6b == io_data_addr[6:0] ? _mem_T_22 : mem_107; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1518 = 7'h6c == io_data_addr[6:0] ? _mem_T_22 : mem_108; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1519 = 7'h6d == io_data_addr[6:0] ? _mem_T_22 : mem_109; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1520 = 7'h6e == io_data_addr[6:0] ? _mem_T_22 : mem_110; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1521 = 7'h6f == io_data_addr[6:0] ? _mem_T_22 : mem_111; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1522 = 7'h70 == io_data_addr[6:0] ? _mem_T_22 : mem_112; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1523 = 7'h71 == io_data_addr[6:0] ? _mem_T_22 : mem_113; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1524 = 7'h72 == io_data_addr[6:0] ? _mem_T_22 : mem_114; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1525 = 7'h73 == io_data_addr[6:0] ? _mem_T_22 : mem_115; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1526 = 7'h74 == io_data_addr[6:0] ? _mem_T_22 : mem_116; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1527 = 7'h75 == io_data_addr[6:0] ? _mem_T_22 : mem_117; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1528 = 7'h76 == io_data_addr[6:0] ? _mem_T_22 : mem_118; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1529 = 7'h77 == io_data_addr[6:0] ? _mem_T_22 : mem_119; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1530 = 7'h78 == io_data_addr[6:0] ? _mem_T_22 : mem_120; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1531 = 7'h79 == io_data_addr[6:0] ? _mem_T_22 : mem_121; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1532 = 7'h7a == io_data_addr[6:0] ? _mem_T_22 : mem_122; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1533 = 7'h7b == io_data_addr[6:0] ? _mem_T_22 : mem_123; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1534 = 7'h7c == io_data_addr[6:0] ? _mem_T_22 : mem_124; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1535 = 7'h7d == io_data_addr[6:0] ? _mem_T_22 : mem_125; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1536 = 7'h7e == io_data_addr[6:0] ? _mem_T_22 : mem_126; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire [31:0] _GEN_1537 = 7'h7f == io_data_addr[6:0] ? _mem_T_22 : mem_127; // @[data.scala 80:25 data.scala 80:25 data.scala 18:16]
  wire  _T_23 = 8'hc == io_data_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_1538 = 7'h0 == io_data_addr[6:0] ? io_data_write : mem_0; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1539 = 7'h1 == io_data_addr[6:0] ? io_data_write : mem_1; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1540 = 7'h2 == io_data_addr[6:0] ? io_data_write : mem_2; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1541 = 7'h3 == io_data_addr[6:0] ? io_data_write : mem_3; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1542 = 7'h4 == io_data_addr[6:0] ? io_data_write : mem_4; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1543 = 7'h5 == io_data_addr[6:0] ? io_data_write : mem_5; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1544 = 7'h6 == io_data_addr[6:0] ? io_data_write : mem_6; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1545 = 7'h7 == io_data_addr[6:0] ? io_data_write : mem_7; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1546 = 7'h8 == io_data_addr[6:0] ? io_data_write : mem_8; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1547 = 7'h9 == io_data_addr[6:0] ? io_data_write : mem_9; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1548 = 7'ha == io_data_addr[6:0] ? io_data_write : mem_10; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1549 = 7'hb == io_data_addr[6:0] ? io_data_write : mem_11; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1550 = 7'hc == io_data_addr[6:0] ? io_data_write : mem_12; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1551 = 7'hd == io_data_addr[6:0] ? io_data_write : mem_13; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1552 = 7'he == io_data_addr[6:0] ? io_data_write : mem_14; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1553 = 7'hf == io_data_addr[6:0] ? io_data_write : mem_15; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1554 = 7'h10 == io_data_addr[6:0] ? io_data_write : mem_16; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1555 = 7'h11 == io_data_addr[6:0] ? io_data_write : mem_17; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1556 = 7'h12 == io_data_addr[6:0] ? io_data_write : mem_18; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1557 = 7'h13 == io_data_addr[6:0] ? io_data_write : mem_19; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1558 = 7'h14 == io_data_addr[6:0] ? io_data_write : mem_20; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1559 = 7'h15 == io_data_addr[6:0] ? io_data_write : mem_21; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1560 = 7'h16 == io_data_addr[6:0] ? io_data_write : mem_22; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1561 = 7'h17 == io_data_addr[6:0] ? io_data_write : mem_23; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1562 = 7'h18 == io_data_addr[6:0] ? io_data_write : mem_24; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1563 = 7'h19 == io_data_addr[6:0] ? io_data_write : mem_25; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1564 = 7'h1a == io_data_addr[6:0] ? io_data_write : mem_26; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1565 = 7'h1b == io_data_addr[6:0] ? io_data_write : mem_27; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1566 = 7'h1c == io_data_addr[6:0] ? io_data_write : mem_28; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1567 = 7'h1d == io_data_addr[6:0] ? io_data_write : mem_29; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1568 = 7'h1e == io_data_addr[6:0] ? io_data_write : mem_30; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1569 = 7'h1f == io_data_addr[6:0] ? io_data_write : mem_31; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1570 = 7'h20 == io_data_addr[6:0] ? io_data_write : mem_32; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1571 = 7'h21 == io_data_addr[6:0] ? io_data_write : mem_33; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1572 = 7'h22 == io_data_addr[6:0] ? io_data_write : mem_34; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1573 = 7'h23 == io_data_addr[6:0] ? io_data_write : mem_35; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1574 = 7'h24 == io_data_addr[6:0] ? io_data_write : mem_36; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1575 = 7'h25 == io_data_addr[6:0] ? io_data_write : mem_37; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1576 = 7'h26 == io_data_addr[6:0] ? io_data_write : mem_38; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1577 = 7'h27 == io_data_addr[6:0] ? io_data_write : mem_39; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1578 = 7'h28 == io_data_addr[6:0] ? io_data_write : mem_40; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1579 = 7'h29 == io_data_addr[6:0] ? io_data_write : mem_41; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1580 = 7'h2a == io_data_addr[6:0] ? io_data_write : mem_42; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1581 = 7'h2b == io_data_addr[6:0] ? io_data_write : mem_43; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1582 = 7'h2c == io_data_addr[6:0] ? io_data_write : mem_44; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1583 = 7'h2d == io_data_addr[6:0] ? io_data_write : mem_45; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1584 = 7'h2e == io_data_addr[6:0] ? io_data_write : mem_46; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1585 = 7'h2f == io_data_addr[6:0] ? io_data_write : mem_47; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1586 = 7'h30 == io_data_addr[6:0] ? io_data_write : mem_48; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1587 = 7'h31 == io_data_addr[6:0] ? io_data_write : mem_49; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1588 = 7'h32 == io_data_addr[6:0] ? io_data_write : mem_50; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1589 = 7'h33 == io_data_addr[6:0] ? io_data_write : mem_51; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1590 = 7'h34 == io_data_addr[6:0] ? io_data_write : mem_52; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1591 = 7'h35 == io_data_addr[6:0] ? io_data_write : mem_53; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1592 = 7'h36 == io_data_addr[6:0] ? io_data_write : mem_54; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1593 = 7'h37 == io_data_addr[6:0] ? io_data_write : mem_55; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1594 = 7'h38 == io_data_addr[6:0] ? io_data_write : mem_56; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1595 = 7'h39 == io_data_addr[6:0] ? io_data_write : mem_57; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1596 = 7'h3a == io_data_addr[6:0] ? io_data_write : mem_58; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1597 = 7'h3b == io_data_addr[6:0] ? io_data_write : mem_59; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1598 = 7'h3c == io_data_addr[6:0] ? io_data_write : mem_60; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1599 = 7'h3d == io_data_addr[6:0] ? io_data_write : mem_61; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1600 = 7'h3e == io_data_addr[6:0] ? io_data_write : mem_62; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1601 = 7'h3f == io_data_addr[6:0] ? io_data_write : mem_63; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1602 = 7'h40 == io_data_addr[6:0] ? io_data_write : mem_64; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1603 = 7'h41 == io_data_addr[6:0] ? io_data_write : mem_65; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1604 = 7'h42 == io_data_addr[6:0] ? io_data_write : mem_66; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1605 = 7'h43 == io_data_addr[6:0] ? io_data_write : mem_67; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1606 = 7'h44 == io_data_addr[6:0] ? io_data_write : mem_68; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1607 = 7'h45 == io_data_addr[6:0] ? io_data_write : mem_69; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1608 = 7'h46 == io_data_addr[6:0] ? io_data_write : mem_70; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1609 = 7'h47 == io_data_addr[6:0] ? io_data_write : mem_71; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1610 = 7'h48 == io_data_addr[6:0] ? io_data_write : mem_72; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1611 = 7'h49 == io_data_addr[6:0] ? io_data_write : mem_73; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1612 = 7'h4a == io_data_addr[6:0] ? io_data_write : mem_74; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1613 = 7'h4b == io_data_addr[6:0] ? io_data_write : mem_75; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1614 = 7'h4c == io_data_addr[6:0] ? io_data_write : mem_76; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1615 = 7'h4d == io_data_addr[6:0] ? io_data_write : mem_77; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1616 = 7'h4e == io_data_addr[6:0] ? io_data_write : mem_78; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1617 = 7'h4f == io_data_addr[6:0] ? io_data_write : mem_79; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1618 = 7'h50 == io_data_addr[6:0] ? io_data_write : mem_80; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1619 = 7'h51 == io_data_addr[6:0] ? io_data_write : mem_81; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1620 = 7'h52 == io_data_addr[6:0] ? io_data_write : mem_82; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1621 = 7'h53 == io_data_addr[6:0] ? io_data_write : mem_83; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1622 = 7'h54 == io_data_addr[6:0] ? io_data_write : mem_84; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1623 = 7'h55 == io_data_addr[6:0] ? io_data_write : mem_85; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1624 = 7'h56 == io_data_addr[6:0] ? io_data_write : mem_86; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1625 = 7'h57 == io_data_addr[6:0] ? io_data_write : mem_87; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1626 = 7'h58 == io_data_addr[6:0] ? io_data_write : mem_88; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1627 = 7'h59 == io_data_addr[6:0] ? io_data_write : mem_89; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1628 = 7'h5a == io_data_addr[6:0] ? io_data_write : mem_90; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1629 = 7'h5b == io_data_addr[6:0] ? io_data_write : mem_91; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1630 = 7'h5c == io_data_addr[6:0] ? io_data_write : mem_92; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1631 = 7'h5d == io_data_addr[6:0] ? io_data_write : mem_93; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1632 = 7'h5e == io_data_addr[6:0] ? io_data_write : mem_94; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1633 = 7'h5f == io_data_addr[6:0] ? io_data_write : mem_95; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1634 = 7'h60 == io_data_addr[6:0] ? io_data_write : mem_96; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1635 = 7'h61 == io_data_addr[6:0] ? io_data_write : mem_97; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1636 = 7'h62 == io_data_addr[6:0] ? io_data_write : mem_98; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1637 = 7'h63 == io_data_addr[6:0] ? io_data_write : mem_99; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1638 = 7'h64 == io_data_addr[6:0] ? io_data_write : mem_100; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1639 = 7'h65 == io_data_addr[6:0] ? io_data_write : mem_101; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1640 = 7'h66 == io_data_addr[6:0] ? io_data_write : mem_102; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1641 = 7'h67 == io_data_addr[6:0] ? io_data_write : mem_103; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1642 = 7'h68 == io_data_addr[6:0] ? io_data_write : mem_104; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1643 = 7'h69 == io_data_addr[6:0] ? io_data_write : mem_105; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1644 = 7'h6a == io_data_addr[6:0] ? io_data_write : mem_106; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1645 = 7'h6b == io_data_addr[6:0] ? io_data_write : mem_107; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1646 = 7'h6c == io_data_addr[6:0] ? io_data_write : mem_108; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1647 = 7'h6d == io_data_addr[6:0] ? io_data_write : mem_109; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1648 = 7'h6e == io_data_addr[6:0] ? io_data_write : mem_110; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1649 = 7'h6f == io_data_addr[6:0] ? io_data_write : mem_111; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1650 = 7'h70 == io_data_addr[6:0] ? io_data_write : mem_112; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1651 = 7'h71 == io_data_addr[6:0] ? io_data_write : mem_113; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1652 = 7'h72 == io_data_addr[6:0] ? io_data_write : mem_114; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1653 = 7'h73 == io_data_addr[6:0] ? io_data_write : mem_115; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1654 = 7'h74 == io_data_addr[6:0] ? io_data_write : mem_116; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1655 = 7'h75 == io_data_addr[6:0] ? io_data_write : mem_117; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1656 = 7'h76 == io_data_addr[6:0] ? io_data_write : mem_118; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1657 = 7'h77 == io_data_addr[6:0] ? io_data_write : mem_119; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1658 = 7'h78 == io_data_addr[6:0] ? io_data_write : mem_120; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1659 = 7'h79 == io_data_addr[6:0] ? io_data_write : mem_121; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1660 = 7'h7a == io_data_addr[6:0] ? io_data_write : mem_122; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1661 = 7'h7b == io_data_addr[6:0] ? io_data_write : mem_123; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1662 = 7'h7c == io_data_addr[6:0] ? io_data_write : mem_124; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1663 = 7'h7d == io_data_addr[6:0] ? io_data_write : mem_125; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1664 = 7'h7e == io_data_addr[6:0] ? io_data_write : mem_126; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1665 = 7'h7f == io_data_addr[6:0] ? io_data_write : mem_127; // @[data.scala 84:25 data.scala 84:25 data.scala 18:16]
  wire [31:0] _GEN_1667 = _T_23 ? _GEN_1538 : mem_0; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1668 = _T_23 ? _GEN_1539 : mem_1; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1669 = _T_23 ? _GEN_1540 : mem_2; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1670 = _T_23 ? _GEN_1541 : mem_3; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1671 = _T_23 ? _GEN_1542 : mem_4; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1672 = _T_23 ? _GEN_1543 : mem_5; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1673 = _T_23 ? _GEN_1544 : mem_6; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1674 = _T_23 ? _GEN_1545 : mem_7; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1675 = _T_23 ? _GEN_1546 : mem_8; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1676 = _T_23 ? _GEN_1547 : mem_9; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1677 = _T_23 ? _GEN_1548 : mem_10; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1678 = _T_23 ? _GEN_1549 : mem_11; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1679 = _T_23 ? _GEN_1550 : mem_12; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1680 = _T_23 ? _GEN_1551 : mem_13; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1681 = _T_23 ? _GEN_1552 : mem_14; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1682 = _T_23 ? _GEN_1553 : mem_15; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1683 = _T_23 ? _GEN_1554 : mem_16; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1684 = _T_23 ? _GEN_1555 : mem_17; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1685 = _T_23 ? _GEN_1556 : mem_18; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1686 = _T_23 ? _GEN_1557 : mem_19; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1687 = _T_23 ? _GEN_1558 : mem_20; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1688 = _T_23 ? _GEN_1559 : mem_21; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1689 = _T_23 ? _GEN_1560 : mem_22; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1690 = _T_23 ? _GEN_1561 : mem_23; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1691 = _T_23 ? _GEN_1562 : mem_24; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1692 = _T_23 ? _GEN_1563 : mem_25; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1693 = _T_23 ? _GEN_1564 : mem_26; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1694 = _T_23 ? _GEN_1565 : mem_27; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1695 = _T_23 ? _GEN_1566 : mem_28; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1696 = _T_23 ? _GEN_1567 : mem_29; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1697 = _T_23 ? _GEN_1568 : mem_30; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1698 = _T_23 ? _GEN_1569 : mem_31; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1699 = _T_23 ? _GEN_1570 : mem_32; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1700 = _T_23 ? _GEN_1571 : mem_33; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1701 = _T_23 ? _GEN_1572 : mem_34; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1702 = _T_23 ? _GEN_1573 : mem_35; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1703 = _T_23 ? _GEN_1574 : mem_36; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1704 = _T_23 ? _GEN_1575 : mem_37; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1705 = _T_23 ? _GEN_1576 : mem_38; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1706 = _T_23 ? _GEN_1577 : mem_39; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1707 = _T_23 ? _GEN_1578 : mem_40; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1708 = _T_23 ? _GEN_1579 : mem_41; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1709 = _T_23 ? _GEN_1580 : mem_42; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1710 = _T_23 ? _GEN_1581 : mem_43; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1711 = _T_23 ? _GEN_1582 : mem_44; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1712 = _T_23 ? _GEN_1583 : mem_45; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1713 = _T_23 ? _GEN_1584 : mem_46; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1714 = _T_23 ? _GEN_1585 : mem_47; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1715 = _T_23 ? _GEN_1586 : mem_48; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1716 = _T_23 ? _GEN_1587 : mem_49; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1717 = _T_23 ? _GEN_1588 : mem_50; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1718 = _T_23 ? _GEN_1589 : mem_51; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1719 = _T_23 ? _GEN_1590 : mem_52; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1720 = _T_23 ? _GEN_1591 : mem_53; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1721 = _T_23 ? _GEN_1592 : mem_54; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1722 = _T_23 ? _GEN_1593 : mem_55; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1723 = _T_23 ? _GEN_1594 : mem_56; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1724 = _T_23 ? _GEN_1595 : mem_57; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1725 = _T_23 ? _GEN_1596 : mem_58; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1726 = _T_23 ? _GEN_1597 : mem_59; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1727 = _T_23 ? _GEN_1598 : mem_60; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1728 = _T_23 ? _GEN_1599 : mem_61; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1729 = _T_23 ? _GEN_1600 : mem_62; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1730 = _T_23 ? _GEN_1601 : mem_63; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1731 = _T_23 ? _GEN_1602 : mem_64; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1732 = _T_23 ? _GEN_1603 : mem_65; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1733 = _T_23 ? _GEN_1604 : mem_66; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1734 = _T_23 ? _GEN_1605 : mem_67; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1735 = _T_23 ? _GEN_1606 : mem_68; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1736 = _T_23 ? _GEN_1607 : mem_69; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1737 = _T_23 ? _GEN_1608 : mem_70; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1738 = _T_23 ? _GEN_1609 : mem_71; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1739 = _T_23 ? _GEN_1610 : mem_72; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1740 = _T_23 ? _GEN_1611 : mem_73; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1741 = _T_23 ? _GEN_1612 : mem_74; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1742 = _T_23 ? _GEN_1613 : mem_75; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1743 = _T_23 ? _GEN_1614 : mem_76; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1744 = _T_23 ? _GEN_1615 : mem_77; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1745 = _T_23 ? _GEN_1616 : mem_78; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1746 = _T_23 ? _GEN_1617 : mem_79; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1747 = _T_23 ? _GEN_1618 : mem_80; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1748 = _T_23 ? _GEN_1619 : mem_81; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1749 = _T_23 ? _GEN_1620 : mem_82; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1750 = _T_23 ? _GEN_1621 : mem_83; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1751 = _T_23 ? _GEN_1622 : mem_84; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1752 = _T_23 ? _GEN_1623 : mem_85; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1753 = _T_23 ? _GEN_1624 : mem_86; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1754 = _T_23 ? _GEN_1625 : mem_87; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1755 = _T_23 ? _GEN_1626 : mem_88; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1756 = _T_23 ? _GEN_1627 : mem_89; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1757 = _T_23 ? _GEN_1628 : mem_90; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1758 = _T_23 ? _GEN_1629 : mem_91; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1759 = _T_23 ? _GEN_1630 : mem_92; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1760 = _T_23 ? _GEN_1631 : mem_93; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1761 = _T_23 ? _GEN_1632 : mem_94; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1762 = _T_23 ? _GEN_1633 : mem_95; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1763 = _T_23 ? _GEN_1634 : mem_96; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1764 = _T_23 ? _GEN_1635 : mem_97; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1765 = _T_23 ? _GEN_1636 : mem_98; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1766 = _T_23 ? _GEN_1637 : mem_99; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1767 = _T_23 ? _GEN_1638 : mem_100; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1768 = _T_23 ? _GEN_1639 : mem_101; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1769 = _T_23 ? _GEN_1640 : mem_102; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1770 = _T_23 ? _GEN_1641 : mem_103; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1771 = _T_23 ? _GEN_1642 : mem_104; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1772 = _T_23 ? _GEN_1643 : mem_105; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1773 = _T_23 ? _GEN_1644 : mem_106; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1774 = _T_23 ? _GEN_1645 : mem_107; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1775 = _T_23 ? _GEN_1646 : mem_108; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1776 = _T_23 ? _GEN_1647 : mem_109; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1777 = _T_23 ? _GEN_1648 : mem_110; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1778 = _T_23 ? _GEN_1649 : mem_111; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1779 = _T_23 ? _GEN_1650 : mem_112; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1780 = _T_23 ? _GEN_1651 : mem_113; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1781 = _T_23 ? _GEN_1652 : mem_114; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1782 = _T_23 ? _GEN_1653 : mem_115; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1783 = _T_23 ? _GEN_1654 : mem_116; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1784 = _T_23 ? _GEN_1655 : mem_117; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1785 = _T_23 ? _GEN_1656 : mem_118; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1786 = _T_23 ? _GEN_1657 : mem_119; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1787 = _T_23 ? _GEN_1658 : mem_120; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1788 = _T_23 ? _GEN_1659 : mem_121; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1789 = _T_23 ? _GEN_1660 : mem_122; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1790 = _T_23 ? _GEN_1661 : mem_123; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1791 = _T_23 ? _GEN_1662 : mem_124; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1792 = _T_23 ? _GEN_1663 : mem_125; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1793 = _T_23 ? _GEN_1664 : mem_126; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1794 = _T_23 ? _GEN_1665 : mem_127; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_1796 = _T_21 ? _GEN_1410 : _GEN_1667; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1797 = _T_21 ? _GEN_1411 : _GEN_1668; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1798 = _T_21 ? _GEN_1412 : _GEN_1669; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1799 = _T_21 ? _GEN_1413 : _GEN_1670; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1800 = _T_21 ? _GEN_1414 : _GEN_1671; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1801 = _T_21 ? _GEN_1415 : _GEN_1672; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1802 = _T_21 ? _GEN_1416 : _GEN_1673; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1803 = _T_21 ? _GEN_1417 : _GEN_1674; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1804 = _T_21 ? _GEN_1418 : _GEN_1675; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1805 = _T_21 ? _GEN_1419 : _GEN_1676; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1806 = _T_21 ? _GEN_1420 : _GEN_1677; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1807 = _T_21 ? _GEN_1421 : _GEN_1678; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1808 = _T_21 ? _GEN_1422 : _GEN_1679; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1809 = _T_21 ? _GEN_1423 : _GEN_1680; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1810 = _T_21 ? _GEN_1424 : _GEN_1681; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1811 = _T_21 ? _GEN_1425 : _GEN_1682; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1812 = _T_21 ? _GEN_1426 : _GEN_1683; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1813 = _T_21 ? _GEN_1427 : _GEN_1684; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1814 = _T_21 ? _GEN_1428 : _GEN_1685; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1815 = _T_21 ? _GEN_1429 : _GEN_1686; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1816 = _T_21 ? _GEN_1430 : _GEN_1687; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1817 = _T_21 ? _GEN_1431 : _GEN_1688; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1818 = _T_21 ? _GEN_1432 : _GEN_1689; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1819 = _T_21 ? _GEN_1433 : _GEN_1690; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1820 = _T_21 ? _GEN_1434 : _GEN_1691; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1821 = _T_21 ? _GEN_1435 : _GEN_1692; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1822 = _T_21 ? _GEN_1436 : _GEN_1693; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1823 = _T_21 ? _GEN_1437 : _GEN_1694; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1824 = _T_21 ? _GEN_1438 : _GEN_1695; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1825 = _T_21 ? _GEN_1439 : _GEN_1696; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1826 = _T_21 ? _GEN_1440 : _GEN_1697; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1827 = _T_21 ? _GEN_1441 : _GEN_1698; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1828 = _T_21 ? _GEN_1442 : _GEN_1699; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1829 = _T_21 ? _GEN_1443 : _GEN_1700; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1830 = _T_21 ? _GEN_1444 : _GEN_1701; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1831 = _T_21 ? _GEN_1445 : _GEN_1702; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1832 = _T_21 ? _GEN_1446 : _GEN_1703; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1833 = _T_21 ? _GEN_1447 : _GEN_1704; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1834 = _T_21 ? _GEN_1448 : _GEN_1705; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1835 = _T_21 ? _GEN_1449 : _GEN_1706; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1836 = _T_21 ? _GEN_1450 : _GEN_1707; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1837 = _T_21 ? _GEN_1451 : _GEN_1708; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1838 = _T_21 ? _GEN_1452 : _GEN_1709; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1839 = _T_21 ? _GEN_1453 : _GEN_1710; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1840 = _T_21 ? _GEN_1454 : _GEN_1711; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1841 = _T_21 ? _GEN_1455 : _GEN_1712; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1842 = _T_21 ? _GEN_1456 : _GEN_1713; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1843 = _T_21 ? _GEN_1457 : _GEN_1714; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1844 = _T_21 ? _GEN_1458 : _GEN_1715; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1845 = _T_21 ? _GEN_1459 : _GEN_1716; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1846 = _T_21 ? _GEN_1460 : _GEN_1717; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1847 = _T_21 ? _GEN_1461 : _GEN_1718; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1848 = _T_21 ? _GEN_1462 : _GEN_1719; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1849 = _T_21 ? _GEN_1463 : _GEN_1720; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1850 = _T_21 ? _GEN_1464 : _GEN_1721; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1851 = _T_21 ? _GEN_1465 : _GEN_1722; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1852 = _T_21 ? _GEN_1466 : _GEN_1723; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1853 = _T_21 ? _GEN_1467 : _GEN_1724; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1854 = _T_21 ? _GEN_1468 : _GEN_1725; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1855 = _T_21 ? _GEN_1469 : _GEN_1726; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1856 = _T_21 ? _GEN_1470 : _GEN_1727; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1857 = _T_21 ? _GEN_1471 : _GEN_1728; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1858 = _T_21 ? _GEN_1472 : _GEN_1729; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1859 = _T_21 ? _GEN_1473 : _GEN_1730; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1860 = _T_21 ? _GEN_1474 : _GEN_1731; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1861 = _T_21 ? _GEN_1475 : _GEN_1732; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1862 = _T_21 ? _GEN_1476 : _GEN_1733; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1863 = _T_21 ? _GEN_1477 : _GEN_1734; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1864 = _T_21 ? _GEN_1478 : _GEN_1735; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1865 = _T_21 ? _GEN_1479 : _GEN_1736; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1866 = _T_21 ? _GEN_1480 : _GEN_1737; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1867 = _T_21 ? _GEN_1481 : _GEN_1738; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1868 = _T_21 ? _GEN_1482 : _GEN_1739; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1869 = _T_21 ? _GEN_1483 : _GEN_1740; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1870 = _T_21 ? _GEN_1484 : _GEN_1741; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1871 = _T_21 ? _GEN_1485 : _GEN_1742; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1872 = _T_21 ? _GEN_1486 : _GEN_1743; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1873 = _T_21 ? _GEN_1487 : _GEN_1744; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1874 = _T_21 ? _GEN_1488 : _GEN_1745; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1875 = _T_21 ? _GEN_1489 : _GEN_1746; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1876 = _T_21 ? _GEN_1490 : _GEN_1747; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1877 = _T_21 ? _GEN_1491 : _GEN_1748; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1878 = _T_21 ? _GEN_1492 : _GEN_1749; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1879 = _T_21 ? _GEN_1493 : _GEN_1750; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1880 = _T_21 ? _GEN_1494 : _GEN_1751; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1881 = _T_21 ? _GEN_1495 : _GEN_1752; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1882 = _T_21 ? _GEN_1496 : _GEN_1753; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1883 = _T_21 ? _GEN_1497 : _GEN_1754; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1884 = _T_21 ? _GEN_1498 : _GEN_1755; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1885 = _T_21 ? _GEN_1499 : _GEN_1756; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1886 = _T_21 ? _GEN_1500 : _GEN_1757; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1887 = _T_21 ? _GEN_1501 : _GEN_1758; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1888 = _T_21 ? _GEN_1502 : _GEN_1759; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1889 = _T_21 ? _GEN_1503 : _GEN_1760; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1890 = _T_21 ? _GEN_1504 : _GEN_1761; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1891 = _T_21 ? _GEN_1505 : _GEN_1762; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1892 = _T_21 ? _GEN_1506 : _GEN_1763; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1893 = _T_21 ? _GEN_1507 : _GEN_1764; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1894 = _T_21 ? _GEN_1508 : _GEN_1765; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1895 = _T_21 ? _GEN_1509 : _GEN_1766; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1896 = _T_21 ? _GEN_1510 : _GEN_1767; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1897 = _T_21 ? _GEN_1511 : _GEN_1768; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1898 = _T_21 ? _GEN_1512 : _GEN_1769; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1899 = _T_21 ? _GEN_1513 : _GEN_1770; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1900 = _T_21 ? _GEN_1514 : _GEN_1771; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1901 = _T_21 ? _GEN_1515 : _GEN_1772; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1902 = _T_21 ? _GEN_1516 : _GEN_1773; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1903 = _T_21 ? _GEN_1517 : _GEN_1774; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1904 = _T_21 ? _GEN_1518 : _GEN_1775; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1905 = _T_21 ? _GEN_1519 : _GEN_1776; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1906 = _T_21 ? _GEN_1520 : _GEN_1777; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1907 = _T_21 ? _GEN_1521 : _GEN_1778; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1908 = _T_21 ? _GEN_1522 : _GEN_1779; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1909 = _T_21 ? _GEN_1523 : _GEN_1780; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1910 = _T_21 ? _GEN_1524 : _GEN_1781; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1911 = _T_21 ? _GEN_1525 : _GEN_1782; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1912 = _T_21 ? _GEN_1526 : _GEN_1783; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1913 = _T_21 ? _GEN_1527 : _GEN_1784; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1914 = _T_21 ? _GEN_1528 : _GEN_1785; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1915 = _T_21 ? _GEN_1529 : _GEN_1786; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1916 = _T_21 ? _GEN_1530 : _GEN_1787; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1917 = _T_21 ? _GEN_1531 : _GEN_1788; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1918 = _T_21 ? _GEN_1532 : _GEN_1789; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1919 = _T_21 ? _GEN_1533 : _GEN_1790; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1920 = _T_21 ? _GEN_1534 : _GEN_1791; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1921 = _T_21 ? _GEN_1535 : _GEN_1792; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1922 = _T_21 ? _GEN_1536 : _GEN_1793; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1923 = _T_21 ? _GEN_1537 : _GEN_1794; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1925 = _T_19 ? _GEN_1282 : _GEN_1796; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1926 = _T_19 ? _GEN_1283 : _GEN_1797; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1927 = _T_19 ? _GEN_1284 : _GEN_1798; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1928 = _T_19 ? _GEN_1285 : _GEN_1799; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1929 = _T_19 ? _GEN_1286 : _GEN_1800; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1930 = _T_19 ? _GEN_1287 : _GEN_1801; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1931 = _T_19 ? _GEN_1288 : _GEN_1802; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1932 = _T_19 ? _GEN_1289 : _GEN_1803; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1933 = _T_19 ? _GEN_1290 : _GEN_1804; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1934 = _T_19 ? _GEN_1291 : _GEN_1805; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1935 = _T_19 ? _GEN_1292 : _GEN_1806; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1936 = _T_19 ? _GEN_1293 : _GEN_1807; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1937 = _T_19 ? _GEN_1294 : _GEN_1808; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1938 = _T_19 ? _GEN_1295 : _GEN_1809; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1939 = _T_19 ? _GEN_1296 : _GEN_1810; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1940 = _T_19 ? _GEN_1297 : _GEN_1811; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1941 = _T_19 ? _GEN_1298 : _GEN_1812; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1942 = _T_19 ? _GEN_1299 : _GEN_1813; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1943 = _T_19 ? _GEN_1300 : _GEN_1814; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1944 = _T_19 ? _GEN_1301 : _GEN_1815; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1945 = _T_19 ? _GEN_1302 : _GEN_1816; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1946 = _T_19 ? _GEN_1303 : _GEN_1817; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1947 = _T_19 ? _GEN_1304 : _GEN_1818; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1948 = _T_19 ? _GEN_1305 : _GEN_1819; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1949 = _T_19 ? _GEN_1306 : _GEN_1820; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1950 = _T_19 ? _GEN_1307 : _GEN_1821; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1951 = _T_19 ? _GEN_1308 : _GEN_1822; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1952 = _T_19 ? _GEN_1309 : _GEN_1823; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1953 = _T_19 ? _GEN_1310 : _GEN_1824; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1954 = _T_19 ? _GEN_1311 : _GEN_1825; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1955 = _T_19 ? _GEN_1312 : _GEN_1826; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1956 = _T_19 ? _GEN_1313 : _GEN_1827; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1957 = _T_19 ? _GEN_1314 : _GEN_1828; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1958 = _T_19 ? _GEN_1315 : _GEN_1829; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1959 = _T_19 ? _GEN_1316 : _GEN_1830; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1960 = _T_19 ? _GEN_1317 : _GEN_1831; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1961 = _T_19 ? _GEN_1318 : _GEN_1832; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1962 = _T_19 ? _GEN_1319 : _GEN_1833; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1963 = _T_19 ? _GEN_1320 : _GEN_1834; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1964 = _T_19 ? _GEN_1321 : _GEN_1835; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1965 = _T_19 ? _GEN_1322 : _GEN_1836; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1966 = _T_19 ? _GEN_1323 : _GEN_1837; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1967 = _T_19 ? _GEN_1324 : _GEN_1838; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1968 = _T_19 ? _GEN_1325 : _GEN_1839; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1969 = _T_19 ? _GEN_1326 : _GEN_1840; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1970 = _T_19 ? _GEN_1327 : _GEN_1841; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1971 = _T_19 ? _GEN_1328 : _GEN_1842; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1972 = _T_19 ? _GEN_1329 : _GEN_1843; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1973 = _T_19 ? _GEN_1330 : _GEN_1844; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1974 = _T_19 ? _GEN_1331 : _GEN_1845; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1975 = _T_19 ? _GEN_1332 : _GEN_1846; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1976 = _T_19 ? _GEN_1333 : _GEN_1847; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1977 = _T_19 ? _GEN_1334 : _GEN_1848; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1978 = _T_19 ? _GEN_1335 : _GEN_1849; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1979 = _T_19 ? _GEN_1336 : _GEN_1850; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1980 = _T_19 ? _GEN_1337 : _GEN_1851; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1981 = _T_19 ? _GEN_1338 : _GEN_1852; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1982 = _T_19 ? _GEN_1339 : _GEN_1853; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1983 = _T_19 ? _GEN_1340 : _GEN_1854; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1984 = _T_19 ? _GEN_1341 : _GEN_1855; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1985 = _T_19 ? _GEN_1342 : _GEN_1856; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1986 = _T_19 ? _GEN_1343 : _GEN_1857; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1987 = _T_19 ? _GEN_1344 : _GEN_1858; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1988 = _T_19 ? _GEN_1345 : _GEN_1859; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1989 = _T_19 ? _GEN_1346 : _GEN_1860; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1990 = _T_19 ? _GEN_1347 : _GEN_1861; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1991 = _T_19 ? _GEN_1348 : _GEN_1862; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1992 = _T_19 ? _GEN_1349 : _GEN_1863; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1993 = _T_19 ? _GEN_1350 : _GEN_1864; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1994 = _T_19 ? _GEN_1351 : _GEN_1865; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1995 = _T_19 ? _GEN_1352 : _GEN_1866; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1996 = _T_19 ? _GEN_1353 : _GEN_1867; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1997 = _T_19 ? _GEN_1354 : _GEN_1868; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1998 = _T_19 ? _GEN_1355 : _GEN_1869; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1999 = _T_19 ? _GEN_1356 : _GEN_1870; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2000 = _T_19 ? _GEN_1357 : _GEN_1871; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2001 = _T_19 ? _GEN_1358 : _GEN_1872; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2002 = _T_19 ? _GEN_1359 : _GEN_1873; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2003 = _T_19 ? _GEN_1360 : _GEN_1874; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2004 = _T_19 ? _GEN_1361 : _GEN_1875; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2005 = _T_19 ? _GEN_1362 : _GEN_1876; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2006 = _T_19 ? _GEN_1363 : _GEN_1877; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2007 = _T_19 ? _GEN_1364 : _GEN_1878; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2008 = _T_19 ? _GEN_1365 : _GEN_1879; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2009 = _T_19 ? _GEN_1366 : _GEN_1880; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2010 = _T_19 ? _GEN_1367 : _GEN_1881; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2011 = _T_19 ? _GEN_1368 : _GEN_1882; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2012 = _T_19 ? _GEN_1369 : _GEN_1883; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2013 = _T_19 ? _GEN_1370 : _GEN_1884; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2014 = _T_19 ? _GEN_1371 : _GEN_1885; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2015 = _T_19 ? _GEN_1372 : _GEN_1886; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2016 = _T_19 ? _GEN_1373 : _GEN_1887; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2017 = _T_19 ? _GEN_1374 : _GEN_1888; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2018 = _T_19 ? _GEN_1375 : _GEN_1889; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2019 = _T_19 ? _GEN_1376 : _GEN_1890; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2020 = _T_19 ? _GEN_1377 : _GEN_1891; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2021 = _T_19 ? _GEN_1378 : _GEN_1892; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2022 = _T_19 ? _GEN_1379 : _GEN_1893; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2023 = _T_19 ? _GEN_1380 : _GEN_1894; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2024 = _T_19 ? _GEN_1381 : _GEN_1895; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2025 = _T_19 ? _GEN_1382 : _GEN_1896; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2026 = _T_19 ? _GEN_1383 : _GEN_1897; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2027 = _T_19 ? _GEN_1384 : _GEN_1898; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2028 = _T_19 ? _GEN_1385 : _GEN_1899; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2029 = _T_19 ? _GEN_1386 : _GEN_1900; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2030 = _T_19 ? _GEN_1387 : _GEN_1901; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2031 = _T_19 ? _GEN_1388 : _GEN_1902; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2032 = _T_19 ? _GEN_1389 : _GEN_1903; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2033 = _T_19 ? _GEN_1390 : _GEN_1904; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2034 = _T_19 ? _GEN_1391 : _GEN_1905; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2035 = _T_19 ? _GEN_1392 : _GEN_1906; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2036 = _T_19 ? _GEN_1393 : _GEN_1907; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2037 = _T_19 ? _GEN_1394 : _GEN_1908; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2038 = _T_19 ? _GEN_1395 : _GEN_1909; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2039 = _T_19 ? _GEN_1396 : _GEN_1910; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2040 = _T_19 ? _GEN_1397 : _GEN_1911; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2041 = _T_19 ? _GEN_1398 : _GEN_1912; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2042 = _T_19 ? _GEN_1399 : _GEN_1913; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2043 = _T_19 ? _GEN_1400 : _GEN_1914; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2044 = _T_19 ? _GEN_1401 : _GEN_1915; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2045 = _T_19 ? _GEN_1402 : _GEN_1916; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2046 = _T_19 ? _GEN_1403 : _GEN_1917; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2047 = _T_19 ? _GEN_1404 : _GEN_1918; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2048 = _T_19 ? _GEN_1405 : _GEN_1919; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2049 = _T_19 ? _GEN_1406 : _GEN_1920; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2050 = _T_19 ? _GEN_1407 : _GEN_1921; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2051 = _T_19 ? _GEN_1408 : _GEN_1922; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2052 = _T_19 ? _GEN_1409 : _GEN_1923; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2054 = _T_18 ? mem_0 : _GEN_1925; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2055 = _T_18 ? mem_1 : _GEN_1926; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2056 = _T_18 ? mem_2 : _GEN_1927; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2057 = _T_18 ? mem_3 : _GEN_1928; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2058 = _T_18 ? mem_4 : _GEN_1929; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2059 = _T_18 ? mem_5 : _GEN_1930; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2060 = _T_18 ? mem_6 : _GEN_1931; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2061 = _T_18 ? mem_7 : _GEN_1932; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2062 = _T_18 ? mem_8 : _GEN_1933; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2063 = _T_18 ? mem_9 : _GEN_1934; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2064 = _T_18 ? mem_10 : _GEN_1935; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2065 = _T_18 ? mem_11 : _GEN_1936; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2066 = _T_18 ? mem_12 : _GEN_1937; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2067 = _T_18 ? mem_13 : _GEN_1938; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2068 = _T_18 ? mem_14 : _GEN_1939; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2069 = _T_18 ? mem_15 : _GEN_1940; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2070 = _T_18 ? mem_16 : _GEN_1941; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2071 = _T_18 ? mem_17 : _GEN_1942; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2072 = _T_18 ? mem_18 : _GEN_1943; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2073 = _T_18 ? mem_19 : _GEN_1944; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2074 = _T_18 ? mem_20 : _GEN_1945; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2075 = _T_18 ? mem_21 : _GEN_1946; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2076 = _T_18 ? mem_22 : _GEN_1947; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2077 = _T_18 ? mem_23 : _GEN_1948; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2078 = _T_18 ? mem_24 : _GEN_1949; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2079 = _T_18 ? mem_25 : _GEN_1950; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2080 = _T_18 ? mem_26 : _GEN_1951; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2081 = _T_18 ? mem_27 : _GEN_1952; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2082 = _T_18 ? mem_28 : _GEN_1953; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2083 = _T_18 ? mem_29 : _GEN_1954; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2084 = _T_18 ? mem_30 : _GEN_1955; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2085 = _T_18 ? mem_31 : _GEN_1956; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2086 = _T_18 ? mem_32 : _GEN_1957; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2087 = _T_18 ? mem_33 : _GEN_1958; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2088 = _T_18 ? mem_34 : _GEN_1959; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2089 = _T_18 ? mem_35 : _GEN_1960; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2090 = _T_18 ? mem_36 : _GEN_1961; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2091 = _T_18 ? mem_37 : _GEN_1962; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2092 = _T_18 ? mem_38 : _GEN_1963; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2093 = _T_18 ? mem_39 : _GEN_1964; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2094 = _T_18 ? mem_40 : _GEN_1965; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2095 = _T_18 ? mem_41 : _GEN_1966; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2096 = _T_18 ? mem_42 : _GEN_1967; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2097 = _T_18 ? mem_43 : _GEN_1968; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2098 = _T_18 ? mem_44 : _GEN_1969; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2099 = _T_18 ? mem_45 : _GEN_1970; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2100 = _T_18 ? mem_46 : _GEN_1971; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2101 = _T_18 ? mem_47 : _GEN_1972; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2102 = _T_18 ? mem_48 : _GEN_1973; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2103 = _T_18 ? mem_49 : _GEN_1974; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2104 = _T_18 ? mem_50 : _GEN_1975; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2105 = _T_18 ? mem_51 : _GEN_1976; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2106 = _T_18 ? mem_52 : _GEN_1977; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2107 = _T_18 ? mem_53 : _GEN_1978; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2108 = _T_18 ? mem_54 : _GEN_1979; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2109 = _T_18 ? mem_55 : _GEN_1980; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2110 = _T_18 ? mem_56 : _GEN_1981; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2111 = _T_18 ? mem_57 : _GEN_1982; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2112 = _T_18 ? mem_58 : _GEN_1983; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2113 = _T_18 ? mem_59 : _GEN_1984; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2114 = _T_18 ? mem_60 : _GEN_1985; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2115 = _T_18 ? mem_61 : _GEN_1986; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2116 = _T_18 ? mem_62 : _GEN_1987; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2117 = _T_18 ? mem_63 : _GEN_1988; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2118 = _T_18 ? mem_64 : _GEN_1989; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2119 = _T_18 ? mem_65 : _GEN_1990; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2120 = _T_18 ? mem_66 : _GEN_1991; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2121 = _T_18 ? mem_67 : _GEN_1992; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2122 = _T_18 ? mem_68 : _GEN_1993; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2123 = _T_18 ? mem_69 : _GEN_1994; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2124 = _T_18 ? mem_70 : _GEN_1995; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2125 = _T_18 ? mem_71 : _GEN_1996; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2126 = _T_18 ? mem_72 : _GEN_1997; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2127 = _T_18 ? mem_73 : _GEN_1998; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2128 = _T_18 ? mem_74 : _GEN_1999; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2129 = _T_18 ? mem_75 : _GEN_2000; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2130 = _T_18 ? mem_76 : _GEN_2001; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2131 = _T_18 ? mem_77 : _GEN_2002; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2132 = _T_18 ? mem_78 : _GEN_2003; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2133 = _T_18 ? mem_79 : _GEN_2004; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2134 = _T_18 ? mem_80 : _GEN_2005; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2135 = _T_18 ? mem_81 : _GEN_2006; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2136 = _T_18 ? mem_82 : _GEN_2007; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2137 = _T_18 ? mem_83 : _GEN_2008; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2138 = _T_18 ? mem_84 : _GEN_2009; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2139 = _T_18 ? mem_85 : _GEN_2010; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2140 = _T_18 ? mem_86 : _GEN_2011; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2141 = _T_18 ? mem_87 : _GEN_2012; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2142 = _T_18 ? mem_88 : _GEN_2013; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2143 = _T_18 ? mem_89 : _GEN_2014; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2144 = _T_18 ? mem_90 : _GEN_2015; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2145 = _T_18 ? mem_91 : _GEN_2016; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2146 = _T_18 ? mem_92 : _GEN_2017; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2147 = _T_18 ? mem_93 : _GEN_2018; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2148 = _T_18 ? mem_94 : _GEN_2019; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2149 = _T_18 ? mem_95 : _GEN_2020; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2150 = _T_18 ? mem_96 : _GEN_2021; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2151 = _T_18 ? mem_97 : _GEN_2022; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2152 = _T_18 ? mem_98 : _GEN_2023; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2153 = _T_18 ? mem_99 : _GEN_2024; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2154 = _T_18 ? mem_100 : _GEN_2025; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2155 = _T_18 ? mem_101 : _GEN_2026; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2156 = _T_18 ? mem_102 : _GEN_2027; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2157 = _T_18 ? mem_103 : _GEN_2028; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2158 = _T_18 ? mem_104 : _GEN_2029; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2159 = _T_18 ? mem_105 : _GEN_2030; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2160 = _T_18 ? mem_106 : _GEN_2031; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2161 = _T_18 ? mem_107 : _GEN_2032; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2162 = _T_18 ? mem_108 : _GEN_2033; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2163 = _T_18 ? mem_109 : _GEN_2034; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2164 = _T_18 ? mem_110 : _GEN_2035; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2165 = _T_18 ? mem_111 : _GEN_2036; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2166 = _T_18 ? mem_112 : _GEN_2037; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2167 = _T_18 ? mem_113 : _GEN_2038; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2168 = _T_18 ? mem_114 : _GEN_2039; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2169 = _T_18 ? mem_115 : _GEN_2040; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2170 = _T_18 ? mem_116 : _GEN_2041; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2171 = _T_18 ? mem_117 : _GEN_2042; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2172 = _T_18 ? mem_118 : _GEN_2043; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2173 = _T_18 ? mem_119 : _GEN_2044; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2174 = _T_18 ? mem_120 : _GEN_2045; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2175 = _T_18 ? mem_121 : _GEN_2046; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2176 = _T_18 ? mem_122 : _GEN_2047; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2177 = _T_18 ? mem_123 : _GEN_2048; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2178 = _T_18 ? mem_124 : _GEN_2049; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2179 = _T_18 ? mem_125 : _GEN_2050; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2180 = _T_18 ? mem_126 : _GEN_2051; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2181 = _T_18 ? mem_127 : _GEN_2052; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2182 = _T_17 ? _GEN_127 : 32'h0; // @[Conditional.scala 39:67 data.scala 69:20]
  wire [31:0] _GEN_2183 = _T_17 ? mem_0 : _GEN_2054; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2184 = _T_17 ? mem_1 : _GEN_2055; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2185 = _T_17 ? mem_2 : _GEN_2056; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2186 = _T_17 ? mem_3 : _GEN_2057; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2187 = _T_17 ? mem_4 : _GEN_2058; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2188 = _T_17 ? mem_5 : _GEN_2059; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2189 = _T_17 ? mem_6 : _GEN_2060; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2190 = _T_17 ? mem_7 : _GEN_2061; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2191 = _T_17 ? mem_8 : _GEN_2062; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2192 = _T_17 ? mem_9 : _GEN_2063; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2193 = _T_17 ? mem_10 : _GEN_2064; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2194 = _T_17 ? mem_11 : _GEN_2065; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2195 = _T_17 ? mem_12 : _GEN_2066; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2196 = _T_17 ? mem_13 : _GEN_2067; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2197 = _T_17 ? mem_14 : _GEN_2068; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2198 = _T_17 ? mem_15 : _GEN_2069; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2199 = _T_17 ? mem_16 : _GEN_2070; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2200 = _T_17 ? mem_17 : _GEN_2071; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2201 = _T_17 ? mem_18 : _GEN_2072; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2202 = _T_17 ? mem_19 : _GEN_2073; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2203 = _T_17 ? mem_20 : _GEN_2074; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2204 = _T_17 ? mem_21 : _GEN_2075; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2205 = _T_17 ? mem_22 : _GEN_2076; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2206 = _T_17 ? mem_23 : _GEN_2077; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2207 = _T_17 ? mem_24 : _GEN_2078; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2208 = _T_17 ? mem_25 : _GEN_2079; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2209 = _T_17 ? mem_26 : _GEN_2080; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2210 = _T_17 ? mem_27 : _GEN_2081; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2211 = _T_17 ? mem_28 : _GEN_2082; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2212 = _T_17 ? mem_29 : _GEN_2083; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2213 = _T_17 ? mem_30 : _GEN_2084; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2214 = _T_17 ? mem_31 : _GEN_2085; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2215 = _T_17 ? mem_32 : _GEN_2086; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2216 = _T_17 ? mem_33 : _GEN_2087; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2217 = _T_17 ? mem_34 : _GEN_2088; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2218 = _T_17 ? mem_35 : _GEN_2089; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2219 = _T_17 ? mem_36 : _GEN_2090; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2220 = _T_17 ? mem_37 : _GEN_2091; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2221 = _T_17 ? mem_38 : _GEN_2092; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2222 = _T_17 ? mem_39 : _GEN_2093; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2223 = _T_17 ? mem_40 : _GEN_2094; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2224 = _T_17 ? mem_41 : _GEN_2095; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2225 = _T_17 ? mem_42 : _GEN_2096; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2226 = _T_17 ? mem_43 : _GEN_2097; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2227 = _T_17 ? mem_44 : _GEN_2098; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2228 = _T_17 ? mem_45 : _GEN_2099; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2229 = _T_17 ? mem_46 : _GEN_2100; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2230 = _T_17 ? mem_47 : _GEN_2101; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2231 = _T_17 ? mem_48 : _GEN_2102; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2232 = _T_17 ? mem_49 : _GEN_2103; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2233 = _T_17 ? mem_50 : _GEN_2104; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2234 = _T_17 ? mem_51 : _GEN_2105; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2235 = _T_17 ? mem_52 : _GEN_2106; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2236 = _T_17 ? mem_53 : _GEN_2107; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2237 = _T_17 ? mem_54 : _GEN_2108; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2238 = _T_17 ? mem_55 : _GEN_2109; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2239 = _T_17 ? mem_56 : _GEN_2110; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2240 = _T_17 ? mem_57 : _GEN_2111; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2241 = _T_17 ? mem_58 : _GEN_2112; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2242 = _T_17 ? mem_59 : _GEN_2113; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2243 = _T_17 ? mem_60 : _GEN_2114; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2244 = _T_17 ? mem_61 : _GEN_2115; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2245 = _T_17 ? mem_62 : _GEN_2116; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2246 = _T_17 ? mem_63 : _GEN_2117; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2247 = _T_17 ? mem_64 : _GEN_2118; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2248 = _T_17 ? mem_65 : _GEN_2119; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2249 = _T_17 ? mem_66 : _GEN_2120; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2250 = _T_17 ? mem_67 : _GEN_2121; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2251 = _T_17 ? mem_68 : _GEN_2122; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2252 = _T_17 ? mem_69 : _GEN_2123; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2253 = _T_17 ? mem_70 : _GEN_2124; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2254 = _T_17 ? mem_71 : _GEN_2125; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2255 = _T_17 ? mem_72 : _GEN_2126; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2256 = _T_17 ? mem_73 : _GEN_2127; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2257 = _T_17 ? mem_74 : _GEN_2128; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2258 = _T_17 ? mem_75 : _GEN_2129; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2259 = _T_17 ? mem_76 : _GEN_2130; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2260 = _T_17 ? mem_77 : _GEN_2131; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2261 = _T_17 ? mem_78 : _GEN_2132; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2262 = _T_17 ? mem_79 : _GEN_2133; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2263 = _T_17 ? mem_80 : _GEN_2134; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2264 = _T_17 ? mem_81 : _GEN_2135; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2265 = _T_17 ? mem_82 : _GEN_2136; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2266 = _T_17 ? mem_83 : _GEN_2137; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2267 = _T_17 ? mem_84 : _GEN_2138; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2268 = _T_17 ? mem_85 : _GEN_2139; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2269 = _T_17 ? mem_86 : _GEN_2140; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2270 = _T_17 ? mem_87 : _GEN_2141; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2271 = _T_17 ? mem_88 : _GEN_2142; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2272 = _T_17 ? mem_89 : _GEN_2143; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2273 = _T_17 ? mem_90 : _GEN_2144; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2274 = _T_17 ? mem_91 : _GEN_2145; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2275 = _T_17 ? mem_92 : _GEN_2146; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2276 = _T_17 ? mem_93 : _GEN_2147; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2277 = _T_17 ? mem_94 : _GEN_2148; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2278 = _T_17 ? mem_95 : _GEN_2149; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2279 = _T_17 ? mem_96 : _GEN_2150; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2280 = _T_17 ? mem_97 : _GEN_2151; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2281 = _T_17 ? mem_98 : _GEN_2152; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2282 = _T_17 ? mem_99 : _GEN_2153; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2283 = _T_17 ? mem_100 : _GEN_2154; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2284 = _T_17 ? mem_101 : _GEN_2155; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2285 = _T_17 ? mem_102 : _GEN_2156; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2286 = _T_17 ? mem_103 : _GEN_2157; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2287 = _T_17 ? mem_104 : _GEN_2158; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2288 = _T_17 ? mem_105 : _GEN_2159; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2289 = _T_17 ? mem_106 : _GEN_2160; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2290 = _T_17 ? mem_107 : _GEN_2161; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2291 = _T_17 ? mem_108 : _GEN_2162; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2292 = _T_17 ? mem_109 : _GEN_2163; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2293 = _T_17 ? mem_110 : _GEN_2164; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2294 = _T_17 ? mem_111 : _GEN_2165; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2295 = _T_17 ? mem_112 : _GEN_2166; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2296 = _T_17 ? mem_113 : _GEN_2167; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2297 = _T_17 ? mem_114 : _GEN_2168; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2298 = _T_17 ? mem_115 : _GEN_2169; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2299 = _T_17 ? mem_116 : _GEN_2170; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2300 = _T_17 ? mem_117 : _GEN_2171; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2301 = _T_17 ? mem_118 : _GEN_2172; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2302 = _T_17 ? mem_119 : _GEN_2173; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2303 = _T_17 ? mem_120 : _GEN_2174; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2304 = _T_17 ? mem_121 : _GEN_2175; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2305 = _T_17 ? mem_122 : _GEN_2176; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2306 = _T_17 ? mem_123 : _GEN_2177; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2307 = _T_17 ? mem_124 : _GEN_2178; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2308 = _T_17 ? mem_125 : _GEN_2179; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2309 = _T_17 ? mem_126 : _GEN_2180; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2310 = _T_17 ? mem_127 : _GEN_2181; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2311 = _T_16 ? _io_data_read_T_18 : _GEN_2182; // @[Conditional.scala 39:67 data.scala 66:20]
  wire [31:0] _GEN_2312 = _T_16 ? mem_0 : _GEN_2183; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2313 = _T_16 ? mem_1 : _GEN_2184; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2314 = _T_16 ? mem_2 : _GEN_2185; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2315 = _T_16 ? mem_3 : _GEN_2186; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2316 = _T_16 ? mem_4 : _GEN_2187; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2317 = _T_16 ? mem_5 : _GEN_2188; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2318 = _T_16 ? mem_6 : _GEN_2189; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2319 = _T_16 ? mem_7 : _GEN_2190; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2320 = _T_16 ? mem_8 : _GEN_2191; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2321 = _T_16 ? mem_9 : _GEN_2192; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2322 = _T_16 ? mem_10 : _GEN_2193; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2323 = _T_16 ? mem_11 : _GEN_2194; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2324 = _T_16 ? mem_12 : _GEN_2195; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2325 = _T_16 ? mem_13 : _GEN_2196; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2326 = _T_16 ? mem_14 : _GEN_2197; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2327 = _T_16 ? mem_15 : _GEN_2198; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2328 = _T_16 ? mem_16 : _GEN_2199; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2329 = _T_16 ? mem_17 : _GEN_2200; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2330 = _T_16 ? mem_18 : _GEN_2201; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2331 = _T_16 ? mem_19 : _GEN_2202; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2332 = _T_16 ? mem_20 : _GEN_2203; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2333 = _T_16 ? mem_21 : _GEN_2204; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2334 = _T_16 ? mem_22 : _GEN_2205; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2335 = _T_16 ? mem_23 : _GEN_2206; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2336 = _T_16 ? mem_24 : _GEN_2207; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2337 = _T_16 ? mem_25 : _GEN_2208; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2338 = _T_16 ? mem_26 : _GEN_2209; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2339 = _T_16 ? mem_27 : _GEN_2210; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2340 = _T_16 ? mem_28 : _GEN_2211; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2341 = _T_16 ? mem_29 : _GEN_2212; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2342 = _T_16 ? mem_30 : _GEN_2213; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2343 = _T_16 ? mem_31 : _GEN_2214; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2344 = _T_16 ? mem_32 : _GEN_2215; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2345 = _T_16 ? mem_33 : _GEN_2216; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2346 = _T_16 ? mem_34 : _GEN_2217; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2347 = _T_16 ? mem_35 : _GEN_2218; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2348 = _T_16 ? mem_36 : _GEN_2219; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2349 = _T_16 ? mem_37 : _GEN_2220; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2350 = _T_16 ? mem_38 : _GEN_2221; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2351 = _T_16 ? mem_39 : _GEN_2222; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2352 = _T_16 ? mem_40 : _GEN_2223; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2353 = _T_16 ? mem_41 : _GEN_2224; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2354 = _T_16 ? mem_42 : _GEN_2225; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2355 = _T_16 ? mem_43 : _GEN_2226; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2356 = _T_16 ? mem_44 : _GEN_2227; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2357 = _T_16 ? mem_45 : _GEN_2228; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2358 = _T_16 ? mem_46 : _GEN_2229; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2359 = _T_16 ? mem_47 : _GEN_2230; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2360 = _T_16 ? mem_48 : _GEN_2231; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2361 = _T_16 ? mem_49 : _GEN_2232; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2362 = _T_16 ? mem_50 : _GEN_2233; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2363 = _T_16 ? mem_51 : _GEN_2234; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2364 = _T_16 ? mem_52 : _GEN_2235; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2365 = _T_16 ? mem_53 : _GEN_2236; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2366 = _T_16 ? mem_54 : _GEN_2237; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2367 = _T_16 ? mem_55 : _GEN_2238; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2368 = _T_16 ? mem_56 : _GEN_2239; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2369 = _T_16 ? mem_57 : _GEN_2240; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2370 = _T_16 ? mem_58 : _GEN_2241; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2371 = _T_16 ? mem_59 : _GEN_2242; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2372 = _T_16 ? mem_60 : _GEN_2243; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2373 = _T_16 ? mem_61 : _GEN_2244; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2374 = _T_16 ? mem_62 : _GEN_2245; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2375 = _T_16 ? mem_63 : _GEN_2246; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2376 = _T_16 ? mem_64 : _GEN_2247; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2377 = _T_16 ? mem_65 : _GEN_2248; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2378 = _T_16 ? mem_66 : _GEN_2249; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2379 = _T_16 ? mem_67 : _GEN_2250; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2380 = _T_16 ? mem_68 : _GEN_2251; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2381 = _T_16 ? mem_69 : _GEN_2252; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2382 = _T_16 ? mem_70 : _GEN_2253; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2383 = _T_16 ? mem_71 : _GEN_2254; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2384 = _T_16 ? mem_72 : _GEN_2255; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2385 = _T_16 ? mem_73 : _GEN_2256; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2386 = _T_16 ? mem_74 : _GEN_2257; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2387 = _T_16 ? mem_75 : _GEN_2258; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2388 = _T_16 ? mem_76 : _GEN_2259; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2389 = _T_16 ? mem_77 : _GEN_2260; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2390 = _T_16 ? mem_78 : _GEN_2261; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2391 = _T_16 ? mem_79 : _GEN_2262; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2392 = _T_16 ? mem_80 : _GEN_2263; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2393 = _T_16 ? mem_81 : _GEN_2264; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2394 = _T_16 ? mem_82 : _GEN_2265; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2395 = _T_16 ? mem_83 : _GEN_2266; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2396 = _T_16 ? mem_84 : _GEN_2267; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2397 = _T_16 ? mem_85 : _GEN_2268; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2398 = _T_16 ? mem_86 : _GEN_2269; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2399 = _T_16 ? mem_87 : _GEN_2270; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2400 = _T_16 ? mem_88 : _GEN_2271; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2401 = _T_16 ? mem_89 : _GEN_2272; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2402 = _T_16 ? mem_90 : _GEN_2273; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2403 = _T_16 ? mem_91 : _GEN_2274; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2404 = _T_16 ? mem_92 : _GEN_2275; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2405 = _T_16 ? mem_93 : _GEN_2276; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2406 = _T_16 ? mem_94 : _GEN_2277; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2407 = _T_16 ? mem_95 : _GEN_2278; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2408 = _T_16 ? mem_96 : _GEN_2279; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2409 = _T_16 ? mem_97 : _GEN_2280; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2410 = _T_16 ? mem_98 : _GEN_2281; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2411 = _T_16 ? mem_99 : _GEN_2282; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2412 = _T_16 ? mem_100 : _GEN_2283; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2413 = _T_16 ? mem_101 : _GEN_2284; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2414 = _T_16 ? mem_102 : _GEN_2285; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2415 = _T_16 ? mem_103 : _GEN_2286; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2416 = _T_16 ? mem_104 : _GEN_2287; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2417 = _T_16 ? mem_105 : _GEN_2288; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2418 = _T_16 ? mem_106 : _GEN_2289; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2419 = _T_16 ? mem_107 : _GEN_2290; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2420 = _T_16 ? mem_108 : _GEN_2291; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2421 = _T_16 ? mem_109 : _GEN_2292; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2422 = _T_16 ? mem_110 : _GEN_2293; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2423 = _T_16 ? mem_111 : _GEN_2294; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2424 = _T_16 ? mem_112 : _GEN_2295; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2425 = _T_16 ? mem_113 : _GEN_2296; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2426 = _T_16 ? mem_114 : _GEN_2297; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2427 = _T_16 ? mem_115 : _GEN_2298; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2428 = _T_16 ? mem_116 : _GEN_2299; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2429 = _T_16 ? mem_117 : _GEN_2300; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2430 = _T_16 ? mem_118 : _GEN_2301; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2431 = _T_16 ? mem_119 : _GEN_2302; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2432 = _T_16 ? mem_120 : _GEN_2303; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2433 = _T_16 ? mem_121 : _GEN_2304; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2434 = _T_16 ? mem_122 : _GEN_2305; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2435 = _T_16 ? mem_123 : _GEN_2306; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2436 = _T_16 ? mem_124 : _GEN_2307; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2437 = _T_16 ? mem_125 : _GEN_2308; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2438 = _T_16 ? mem_126 : _GEN_2309; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2439 = _T_16 ? mem_127 : _GEN_2310; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2440 = _T_15 ? {{16'd0}, _GEN_127[15:0]} : _GEN_2311; // @[Conditional.scala 39:67 data.scala 63:20]
  wire [31:0] _GEN_2441 = _T_15 ? mem_0 : _GEN_2312; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2442 = _T_15 ? mem_1 : _GEN_2313; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2443 = _T_15 ? mem_2 : _GEN_2314; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2444 = _T_15 ? mem_3 : _GEN_2315; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2445 = _T_15 ? mem_4 : _GEN_2316; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2446 = _T_15 ? mem_5 : _GEN_2317; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2447 = _T_15 ? mem_6 : _GEN_2318; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2448 = _T_15 ? mem_7 : _GEN_2319; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2449 = _T_15 ? mem_8 : _GEN_2320; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2450 = _T_15 ? mem_9 : _GEN_2321; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2451 = _T_15 ? mem_10 : _GEN_2322; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2452 = _T_15 ? mem_11 : _GEN_2323; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2453 = _T_15 ? mem_12 : _GEN_2324; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2454 = _T_15 ? mem_13 : _GEN_2325; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2455 = _T_15 ? mem_14 : _GEN_2326; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2456 = _T_15 ? mem_15 : _GEN_2327; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2457 = _T_15 ? mem_16 : _GEN_2328; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2458 = _T_15 ? mem_17 : _GEN_2329; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2459 = _T_15 ? mem_18 : _GEN_2330; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2460 = _T_15 ? mem_19 : _GEN_2331; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2461 = _T_15 ? mem_20 : _GEN_2332; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2462 = _T_15 ? mem_21 : _GEN_2333; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2463 = _T_15 ? mem_22 : _GEN_2334; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2464 = _T_15 ? mem_23 : _GEN_2335; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2465 = _T_15 ? mem_24 : _GEN_2336; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2466 = _T_15 ? mem_25 : _GEN_2337; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2467 = _T_15 ? mem_26 : _GEN_2338; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2468 = _T_15 ? mem_27 : _GEN_2339; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2469 = _T_15 ? mem_28 : _GEN_2340; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2470 = _T_15 ? mem_29 : _GEN_2341; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2471 = _T_15 ? mem_30 : _GEN_2342; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2472 = _T_15 ? mem_31 : _GEN_2343; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2473 = _T_15 ? mem_32 : _GEN_2344; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2474 = _T_15 ? mem_33 : _GEN_2345; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2475 = _T_15 ? mem_34 : _GEN_2346; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2476 = _T_15 ? mem_35 : _GEN_2347; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2477 = _T_15 ? mem_36 : _GEN_2348; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2478 = _T_15 ? mem_37 : _GEN_2349; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2479 = _T_15 ? mem_38 : _GEN_2350; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2480 = _T_15 ? mem_39 : _GEN_2351; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2481 = _T_15 ? mem_40 : _GEN_2352; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2482 = _T_15 ? mem_41 : _GEN_2353; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2483 = _T_15 ? mem_42 : _GEN_2354; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2484 = _T_15 ? mem_43 : _GEN_2355; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2485 = _T_15 ? mem_44 : _GEN_2356; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2486 = _T_15 ? mem_45 : _GEN_2357; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2487 = _T_15 ? mem_46 : _GEN_2358; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2488 = _T_15 ? mem_47 : _GEN_2359; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2489 = _T_15 ? mem_48 : _GEN_2360; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2490 = _T_15 ? mem_49 : _GEN_2361; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2491 = _T_15 ? mem_50 : _GEN_2362; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2492 = _T_15 ? mem_51 : _GEN_2363; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2493 = _T_15 ? mem_52 : _GEN_2364; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2494 = _T_15 ? mem_53 : _GEN_2365; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2495 = _T_15 ? mem_54 : _GEN_2366; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2496 = _T_15 ? mem_55 : _GEN_2367; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2497 = _T_15 ? mem_56 : _GEN_2368; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2498 = _T_15 ? mem_57 : _GEN_2369; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2499 = _T_15 ? mem_58 : _GEN_2370; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2500 = _T_15 ? mem_59 : _GEN_2371; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2501 = _T_15 ? mem_60 : _GEN_2372; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2502 = _T_15 ? mem_61 : _GEN_2373; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2503 = _T_15 ? mem_62 : _GEN_2374; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2504 = _T_15 ? mem_63 : _GEN_2375; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2505 = _T_15 ? mem_64 : _GEN_2376; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2506 = _T_15 ? mem_65 : _GEN_2377; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2507 = _T_15 ? mem_66 : _GEN_2378; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2508 = _T_15 ? mem_67 : _GEN_2379; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2509 = _T_15 ? mem_68 : _GEN_2380; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2510 = _T_15 ? mem_69 : _GEN_2381; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2511 = _T_15 ? mem_70 : _GEN_2382; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2512 = _T_15 ? mem_71 : _GEN_2383; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2513 = _T_15 ? mem_72 : _GEN_2384; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2514 = _T_15 ? mem_73 : _GEN_2385; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2515 = _T_15 ? mem_74 : _GEN_2386; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2516 = _T_15 ? mem_75 : _GEN_2387; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2517 = _T_15 ? mem_76 : _GEN_2388; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2518 = _T_15 ? mem_77 : _GEN_2389; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2519 = _T_15 ? mem_78 : _GEN_2390; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2520 = _T_15 ? mem_79 : _GEN_2391; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2521 = _T_15 ? mem_80 : _GEN_2392; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2522 = _T_15 ? mem_81 : _GEN_2393; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2523 = _T_15 ? mem_82 : _GEN_2394; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2524 = _T_15 ? mem_83 : _GEN_2395; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2525 = _T_15 ? mem_84 : _GEN_2396; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2526 = _T_15 ? mem_85 : _GEN_2397; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2527 = _T_15 ? mem_86 : _GEN_2398; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2528 = _T_15 ? mem_87 : _GEN_2399; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2529 = _T_15 ? mem_88 : _GEN_2400; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2530 = _T_15 ? mem_89 : _GEN_2401; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2531 = _T_15 ? mem_90 : _GEN_2402; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2532 = _T_15 ? mem_91 : _GEN_2403; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2533 = _T_15 ? mem_92 : _GEN_2404; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2534 = _T_15 ? mem_93 : _GEN_2405; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2535 = _T_15 ? mem_94 : _GEN_2406; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2536 = _T_15 ? mem_95 : _GEN_2407; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2537 = _T_15 ? mem_96 : _GEN_2408; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2538 = _T_15 ? mem_97 : _GEN_2409; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2539 = _T_15 ? mem_98 : _GEN_2410; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2540 = _T_15 ? mem_99 : _GEN_2411; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2541 = _T_15 ? mem_100 : _GEN_2412; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2542 = _T_15 ? mem_101 : _GEN_2413; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2543 = _T_15 ? mem_102 : _GEN_2414; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2544 = _T_15 ? mem_103 : _GEN_2415; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2545 = _T_15 ? mem_104 : _GEN_2416; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2546 = _T_15 ? mem_105 : _GEN_2417; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2547 = _T_15 ? mem_106 : _GEN_2418; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2548 = _T_15 ? mem_107 : _GEN_2419; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2549 = _T_15 ? mem_108 : _GEN_2420; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2550 = _T_15 ? mem_109 : _GEN_2421; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2551 = _T_15 ? mem_110 : _GEN_2422; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2552 = _T_15 ? mem_111 : _GEN_2423; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2553 = _T_15 ? mem_112 : _GEN_2424; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2554 = _T_15 ? mem_113 : _GEN_2425; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2555 = _T_15 ? mem_114 : _GEN_2426; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2556 = _T_15 ? mem_115 : _GEN_2427; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2557 = _T_15 ? mem_116 : _GEN_2428; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2558 = _T_15 ? mem_117 : _GEN_2429; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2559 = _T_15 ? mem_118 : _GEN_2430; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2560 = _T_15 ? mem_119 : _GEN_2431; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2561 = _T_15 ? mem_120 : _GEN_2432; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2562 = _T_15 ? mem_121 : _GEN_2433; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2563 = _T_15 ? mem_122 : _GEN_2434; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2564 = _T_15 ? mem_123 : _GEN_2435; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2565 = _T_15 ? mem_124 : _GEN_2436; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2566 = _T_15 ? mem_125 : _GEN_2437; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2567 = _T_15 ? mem_126 : _GEN_2438; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2568 = _T_15 ? mem_127 : _GEN_2439; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2569 = _T_11 ? _GEN_897 : _GEN_2440; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2570 = _T_11 ? mem_0 : _GEN_2441; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2571 = _T_11 ? mem_1 : _GEN_2442; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2572 = _T_11 ? mem_2 : _GEN_2443; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2573 = _T_11 ? mem_3 : _GEN_2444; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2574 = _T_11 ? mem_4 : _GEN_2445; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2575 = _T_11 ? mem_5 : _GEN_2446; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2576 = _T_11 ? mem_6 : _GEN_2447; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2577 = _T_11 ? mem_7 : _GEN_2448; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2578 = _T_11 ? mem_8 : _GEN_2449; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2579 = _T_11 ? mem_9 : _GEN_2450; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2580 = _T_11 ? mem_10 : _GEN_2451; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2581 = _T_11 ? mem_11 : _GEN_2452; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2582 = _T_11 ? mem_12 : _GEN_2453; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2583 = _T_11 ? mem_13 : _GEN_2454; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2584 = _T_11 ? mem_14 : _GEN_2455; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2585 = _T_11 ? mem_15 : _GEN_2456; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2586 = _T_11 ? mem_16 : _GEN_2457; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2587 = _T_11 ? mem_17 : _GEN_2458; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2588 = _T_11 ? mem_18 : _GEN_2459; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2589 = _T_11 ? mem_19 : _GEN_2460; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2590 = _T_11 ? mem_20 : _GEN_2461; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2591 = _T_11 ? mem_21 : _GEN_2462; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2592 = _T_11 ? mem_22 : _GEN_2463; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2593 = _T_11 ? mem_23 : _GEN_2464; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2594 = _T_11 ? mem_24 : _GEN_2465; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2595 = _T_11 ? mem_25 : _GEN_2466; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2596 = _T_11 ? mem_26 : _GEN_2467; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2597 = _T_11 ? mem_27 : _GEN_2468; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2598 = _T_11 ? mem_28 : _GEN_2469; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2599 = _T_11 ? mem_29 : _GEN_2470; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2600 = _T_11 ? mem_30 : _GEN_2471; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2601 = _T_11 ? mem_31 : _GEN_2472; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2602 = _T_11 ? mem_32 : _GEN_2473; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2603 = _T_11 ? mem_33 : _GEN_2474; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2604 = _T_11 ? mem_34 : _GEN_2475; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2605 = _T_11 ? mem_35 : _GEN_2476; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2606 = _T_11 ? mem_36 : _GEN_2477; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2607 = _T_11 ? mem_37 : _GEN_2478; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2608 = _T_11 ? mem_38 : _GEN_2479; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2609 = _T_11 ? mem_39 : _GEN_2480; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2610 = _T_11 ? mem_40 : _GEN_2481; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2611 = _T_11 ? mem_41 : _GEN_2482; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2612 = _T_11 ? mem_42 : _GEN_2483; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2613 = _T_11 ? mem_43 : _GEN_2484; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2614 = _T_11 ? mem_44 : _GEN_2485; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2615 = _T_11 ? mem_45 : _GEN_2486; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2616 = _T_11 ? mem_46 : _GEN_2487; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2617 = _T_11 ? mem_47 : _GEN_2488; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2618 = _T_11 ? mem_48 : _GEN_2489; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2619 = _T_11 ? mem_49 : _GEN_2490; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2620 = _T_11 ? mem_50 : _GEN_2491; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2621 = _T_11 ? mem_51 : _GEN_2492; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2622 = _T_11 ? mem_52 : _GEN_2493; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2623 = _T_11 ? mem_53 : _GEN_2494; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2624 = _T_11 ? mem_54 : _GEN_2495; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2625 = _T_11 ? mem_55 : _GEN_2496; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2626 = _T_11 ? mem_56 : _GEN_2497; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2627 = _T_11 ? mem_57 : _GEN_2498; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2628 = _T_11 ? mem_58 : _GEN_2499; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2629 = _T_11 ? mem_59 : _GEN_2500; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2630 = _T_11 ? mem_60 : _GEN_2501; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2631 = _T_11 ? mem_61 : _GEN_2502; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2632 = _T_11 ? mem_62 : _GEN_2503; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2633 = _T_11 ? mem_63 : _GEN_2504; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2634 = _T_11 ? mem_64 : _GEN_2505; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2635 = _T_11 ? mem_65 : _GEN_2506; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2636 = _T_11 ? mem_66 : _GEN_2507; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2637 = _T_11 ? mem_67 : _GEN_2508; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2638 = _T_11 ? mem_68 : _GEN_2509; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2639 = _T_11 ? mem_69 : _GEN_2510; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2640 = _T_11 ? mem_70 : _GEN_2511; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2641 = _T_11 ? mem_71 : _GEN_2512; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2642 = _T_11 ? mem_72 : _GEN_2513; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2643 = _T_11 ? mem_73 : _GEN_2514; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2644 = _T_11 ? mem_74 : _GEN_2515; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2645 = _T_11 ? mem_75 : _GEN_2516; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2646 = _T_11 ? mem_76 : _GEN_2517; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2647 = _T_11 ? mem_77 : _GEN_2518; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2648 = _T_11 ? mem_78 : _GEN_2519; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2649 = _T_11 ? mem_79 : _GEN_2520; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2650 = _T_11 ? mem_80 : _GEN_2521; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2651 = _T_11 ? mem_81 : _GEN_2522; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2652 = _T_11 ? mem_82 : _GEN_2523; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2653 = _T_11 ? mem_83 : _GEN_2524; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2654 = _T_11 ? mem_84 : _GEN_2525; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2655 = _T_11 ? mem_85 : _GEN_2526; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2656 = _T_11 ? mem_86 : _GEN_2527; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2657 = _T_11 ? mem_87 : _GEN_2528; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2658 = _T_11 ? mem_88 : _GEN_2529; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2659 = _T_11 ? mem_89 : _GEN_2530; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2660 = _T_11 ? mem_90 : _GEN_2531; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2661 = _T_11 ? mem_91 : _GEN_2532; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2662 = _T_11 ? mem_92 : _GEN_2533; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2663 = _T_11 ? mem_93 : _GEN_2534; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2664 = _T_11 ? mem_94 : _GEN_2535; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2665 = _T_11 ? mem_95 : _GEN_2536; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2666 = _T_11 ? mem_96 : _GEN_2537; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2667 = _T_11 ? mem_97 : _GEN_2538; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2668 = _T_11 ? mem_98 : _GEN_2539; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2669 = _T_11 ? mem_99 : _GEN_2540; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2670 = _T_11 ? mem_100 : _GEN_2541; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2671 = _T_11 ? mem_101 : _GEN_2542; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2672 = _T_11 ? mem_102 : _GEN_2543; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2673 = _T_11 ? mem_103 : _GEN_2544; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2674 = _T_11 ? mem_104 : _GEN_2545; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2675 = _T_11 ? mem_105 : _GEN_2546; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2676 = _T_11 ? mem_106 : _GEN_2547; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2677 = _T_11 ? mem_107 : _GEN_2548; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2678 = _T_11 ? mem_108 : _GEN_2549; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2679 = _T_11 ? mem_109 : _GEN_2550; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2680 = _T_11 ? mem_110 : _GEN_2551; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2681 = _T_11 ? mem_111 : _GEN_2552; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2682 = _T_11 ? mem_112 : _GEN_2553; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2683 = _T_11 ? mem_113 : _GEN_2554; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2684 = _T_11 ? mem_114 : _GEN_2555; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2685 = _T_11 ? mem_115 : _GEN_2556; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2686 = _T_11 ? mem_116 : _GEN_2557; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2687 = _T_11 ? mem_117 : _GEN_2558; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2688 = _T_11 ? mem_118 : _GEN_2559; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2689 = _T_11 ? mem_119 : _GEN_2560; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2690 = _T_11 ? mem_120 : _GEN_2561; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2691 = _T_11 ? mem_121 : _GEN_2562; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2692 = _T_11 ? mem_122 : _GEN_2563; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2693 = _T_11 ? mem_123 : _GEN_2564; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2694 = _T_11 ? mem_124 : _GEN_2565; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2695 = _T_11 ? mem_125 : _GEN_2566; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2696 = _T_11 ? mem_126 : _GEN_2567; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2697 = _T_11 ? mem_127 : _GEN_2568; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2698 = _T_10 ? {{24'd0}, _GEN_127[7:0]} : _GEN_2569; // @[Conditional.scala 39:67 data.scala 52:20]
  wire [31:0] _GEN_2699 = _T_10 ? mem_0 : _GEN_2570; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2700 = _T_10 ? mem_1 : _GEN_2571; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2701 = _T_10 ? mem_2 : _GEN_2572; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2702 = _T_10 ? mem_3 : _GEN_2573; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2703 = _T_10 ? mem_4 : _GEN_2574; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2704 = _T_10 ? mem_5 : _GEN_2575; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2705 = _T_10 ? mem_6 : _GEN_2576; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2706 = _T_10 ? mem_7 : _GEN_2577; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2707 = _T_10 ? mem_8 : _GEN_2578; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2708 = _T_10 ? mem_9 : _GEN_2579; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2709 = _T_10 ? mem_10 : _GEN_2580; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2710 = _T_10 ? mem_11 : _GEN_2581; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2711 = _T_10 ? mem_12 : _GEN_2582; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2712 = _T_10 ? mem_13 : _GEN_2583; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2713 = _T_10 ? mem_14 : _GEN_2584; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2714 = _T_10 ? mem_15 : _GEN_2585; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2715 = _T_10 ? mem_16 : _GEN_2586; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2716 = _T_10 ? mem_17 : _GEN_2587; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2717 = _T_10 ? mem_18 : _GEN_2588; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2718 = _T_10 ? mem_19 : _GEN_2589; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2719 = _T_10 ? mem_20 : _GEN_2590; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2720 = _T_10 ? mem_21 : _GEN_2591; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2721 = _T_10 ? mem_22 : _GEN_2592; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2722 = _T_10 ? mem_23 : _GEN_2593; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2723 = _T_10 ? mem_24 : _GEN_2594; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2724 = _T_10 ? mem_25 : _GEN_2595; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2725 = _T_10 ? mem_26 : _GEN_2596; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2726 = _T_10 ? mem_27 : _GEN_2597; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2727 = _T_10 ? mem_28 : _GEN_2598; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2728 = _T_10 ? mem_29 : _GEN_2599; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2729 = _T_10 ? mem_30 : _GEN_2600; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2730 = _T_10 ? mem_31 : _GEN_2601; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2731 = _T_10 ? mem_32 : _GEN_2602; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2732 = _T_10 ? mem_33 : _GEN_2603; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2733 = _T_10 ? mem_34 : _GEN_2604; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2734 = _T_10 ? mem_35 : _GEN_2605; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2735 = _T_10 ? mem_36 : _GEN_2606; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2736 = _T_10 ? mem_37 : _GEN_2607; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2737 = _T_10 ? mem_38 : _GEN_2608; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2738 = _T_10 ? mem_39 : _GEN_2609; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2739 = _T_10 ? mem_40 : _GEN_2610; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2740 = _T_10 ? mem_41 : _GEN_2611; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2741 = _T_10 ? mem_42 : _GEN_2612; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2742 = _T_10 ? mem_43 : _GEN_2613; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2743 = _T_10 ? mem_44 : _GEN_2614; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2744 = _T_10 ? mem_45 : _GEN_2615; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2745 = _T_10 ? mem_46 : _GEN_2616; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2746 = _T_10 ? mem_47 : _GEN_2617; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2747 = _T_10 ? mem_48 : _GEN_2618; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2748 = _T_10 ? mem_49 : _GEN_2619; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2749 = _T_10 ? mem_50 : _GEN_2620; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2750 = _T_10 ? mem_51 : _GEN_2621; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2751 = _T_10 ? mem_52 : _GEN_2622; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2752 = _T_10 ? mem_53 : _GEN_2623; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2753 = _T_10 ? mem_54 : _GEN_2624; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2754 = _T_10 ? mem_55 : _GEN_2625; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2755 = _T_10 ? mem_56 : _GEN_2626; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2756 = _T_10 ? mem_57 : _GEN_2627; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2757 = _T_10 ? mem_58 : _GEN_2628; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2758 = _T_10 ? mem_59 : _GEN_2629; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2759 = _T_10 ? mem_60 : _GEN_2630; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2760 = _T_10 ? mem_61 : _GEN_2631; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2761 = _T_10 ? mem_62 : _GEN_2632; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2762 = _T_10 ? mem_63 : _GEN_2633; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2763 = _T_10 ? mem_64 : _GEN_2634; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2764 = _T_10 ? mem_65 : _GEN_2635; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2765 = _T_10 ? mem_66 : _GEN_2636; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2766 = _T_10 ? mem_67 : _GEN_2637; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2767 = _T_10 ? mem_68 : _GEN_2638; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2768 = _T_10 ? mem_69 : _GEN_2639; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2769 = _T_10 ? mem_70 : _GEN_2640; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2770 = _T_10 ? mem_71 : _GEN_2641; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2771 = _T_10 ? mem_72 : _GEN_2642; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2772 = _T_10 ? mem_73 : _GEN_2643; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2773 = _T_10 ? mem_74 : _GEN_2644; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2774 = _T_10 ? mem_75 : _GEN_2645; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2775 = _T_10 ? mem_76 : _GEN_2646; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2776 = _T_10 ? mem_77 : _GEN_2647; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2777 = _T_10 ? mem_78 : _GEN_2648; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2778 = _T_10 ? mem_79 : _GEN_2649; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2779 = _T_10 ? mem_80 : _GEN_2650; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2780 = _T_10 ? mem_81 : _GEN_2651; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2781 = _T_10 ? mem_82 : _GEN_2652; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2782 = _T_10 ? mem_83 : _GEN_2653; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2783 = _T_10 ? mem_84 : _GEN_2654; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2784 = _T_10 ? mem_85 : _GEN_2655; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2785 = _T_10 ? mem_86 : _GEN_2656; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2786 = _T_10 ? mem_87 : _GEN_2657; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2787 = _T_10 ? mem_88 : _GEN_2658; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2788 = _T_10 ? mem_89 : _GEN_2659; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2789 = _T_10 ? mem_90 : _GEN_2660; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2790 = _T_10 ? mem_91 : _GEN_2661; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2791 = _T_10 ? mem_92 : _GEN_2662; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2792 = _T_10 ? mem_93 : _GEN_2663; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2793 = _T_10 ? mem_94 : _GEN_2664; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2794 = _T_10 ? mem_95 : _GEN_2665; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2795 = _T_10 ? mem_96 : _GEN_2666; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2796 = _T_10 ? mem_97 : _GEN_2667; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2797 = _T_10 ? mem_98 : _GEN_2668; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2798 = _T_10 ? mem_99 : _GEN_2669; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2799 = _T_10 ? mem_100 : _GEN_2670; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2800 = _T_10 ? mem_101 : _GEN_2671; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2801 = _T_10 ? mem_102 : _GEN_2672; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2802 = _T_10 ? mem_103 : _GEN_2673; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2803 = _T_10 ? mem_104 : _GEN_2674; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2804 = _T_10 ? mem_105 : _GEN_2675; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2805 = _T_10 ? mem_106 : _GEN_2676; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2806 = _T_10 ? mem_107 : _GEN_2677; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2807 = _T_10 ? mem_108 : _GEN_2678; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2808 = _T_10 ? mem_109 : _GEN_2679; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2809 = _T_10 ? mem_110 : _GEN_2680; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2810 = _T_10 ? mem_111 : _GEN_2681; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2811 = _T_10 ? mem_112 : _GEN_2682; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2812 = _T_10 ? mem_113 : _GEN_2683; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2813 = _T_10 ? mem_114 : _GEN_2684; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2814 = _T_10 ? mem_115 : _GEN_2685; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2815 = _T_10 ? mem_116 : _GEN_2686; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2816 = _T_10 ? mem_117 : _GEN_2687; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2817 = _T_10 ? mem_118 : _GEN_2688; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2818 = _T_10 ? mem_119 : _GEN_2689; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2819 = _T_10 ? mem_120 : _GEN_2690; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2820 = _T_10 ? mem_121 : _GEN_2691; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2821 = _T_10 ? mem_122 : _GEN_2692; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2822 = _T_10 ? mem_123 : _GEN_2693; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2823 = _T_10 ? mem_124 : _GEN_2694; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2824 = _T_10 ? mem_125 : _GEN_2695; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2825 = _T_10 ? mem_126 : _GEN_2696; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2826 = _T_10 ? mem_127 : _GEN_2697; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2827 = _T_6 ? _GEN_384 : _GEN_2698; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2828 = _T_6 ? mem_0 : _GEN_2699; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2829 = _T_6 ? mem_1 : _GEN_2700; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2830 = _T_6 ? mem_2 : _GEN_2701; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2831 = _T_6 ? mem_3 : _GEN_2702; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2832 = _T_6 ? mem_4 : _GEN_2703; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2833 = _T_6 ? mem_5 : _GEN_2704; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2834 = _T_6 ? mem_6 : _GEN_2705; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2835 = _T_6 ? mem_7 : _GEN_2706; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2836 = _T_6 ? mem_8 : _GEN_2707; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2837 = _T_6 ? mem_9 : _GEN_2708; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2838 = _T_6 ? mem_10 : _GEN_2709; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2839 = _T_6 ? mem_11 : _GEN_2710; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2840 = _T_6 ? mem_12 : _GEN_2711; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2841 = _T_6 ? mem_13 : _GEN_2712; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2842 = _T_6 ? mem_14 : _GEN_2713; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2843 = _T_6 ? mem_15 : _GEN_2714; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2844 = _T_6 ? mem_16 : _GEN_2715; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2845 = _T_6 ? mem_17 : _GEN_2716; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2846 = _T_6 ? mem_18 : _GEN_2717; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2847 = _T_6 ? mem_19 : _GEN_2718; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2848 = _T_6 ? mem_20 : _GEN_2719; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2849 = _T_6 ? mem_21 : _GEN_2720; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2850 = _T_6 ? mem_22 : _GEN_2721; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2851 = _T_6 ? mem_23 : _GEN_2722; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2852 = _T_6 ? mem_24 : _GEN_2723; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2853 = _T_6 ? mem_25 : _GEN_2724; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2854 = _T_6 ? mem_26 : _GEN_2725; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2855 = _T_6 ? mem_27 : _GEN_2726; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2856 = _T_6 ? mem_28 : _GEN_2727; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2857 = _T_6 ? mem_29 : _GEN_2728; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2858 = _T_6 ? mem_30 : _GEN_2729; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2859 = _T_6 ? mem_31 : _GEN_2730; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2860 = _T_6 ? mem_32 : _GEN_2731; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2861 = _T_6 ? mem_33 : _GEN_2732; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2862 = _T_6 ? mem_34 : _GEN_2733; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2863 = _T_6 ? mem_35 : _GEN_2734; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2864 = _T_6 ? mem_36 : _GEN_2735; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2865 = _T_6 ? mem_37 : _GEN_2736; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2866 = _T_6 ? mem_38 : _GEN_2737; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2867 = _T_6 ? mem_39 : _GEN_2738; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2868 = _T_6 ? mem_40 : _GEN_2739; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2869 = _T_6 ? mem_41 : _GEN_2740; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2870 = _T_6 ? mem_42 : _GEN_2741; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2871 = _T_6 ? mem_43 : _GEN_2742; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2872 = _T_6 ? mem_44 : _GEN_2743; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2873 = _T_6 ? mem_45 : _GEN_2744; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2874 = _T_6 ? mem_46 : _GEN_2745; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2875 = _T_6 ? mem_47 : _GEN_2746; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2876 = _T_6 ? mem_48 : _GEN_2747; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2877 = _T_6 ? mem_49 : _GEN_2748; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2878 = _T_6 ? mem_50 : _GEN_2749; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2879 = _T_6 ? mem_51 : _GEN_2750; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2880 = _T_6 ? mem_52 : _GEN_2751; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2881 = _T_6 ? mem_53 : _GEN_2752; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2882 = _T_6 ? mem_54 : _GEN_2753; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2883 = _T_6 ? mem_55 : _GEN_2754; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2884 = _T_6 ? mem_56 : _GEN_2755; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2885 = _T_6 ? mem_57 : _GEN_2756; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2886 = _T_6 ? mem_58 : _GEN_2757; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2887 = _T_6 ? mem_59 : _GEN_2758; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2888 = _T_6 ? mem_60 : _GEN_2759; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2889 = _T_6 ? mem_61 : _GEN_2760; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2890 = _T_6 ? mem_62 : _GEN_2761; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2891 = _T_6 ? mem_63 : _GEN_2762; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2892 = _T_6 ? mem_64 : _GEN_2763; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2893 = _T_6 ? mem_65 : _GEN_2764; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2894 = _T_6 ? mem_66 : _GEN_2765; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2895 = _T_6 ? mem_67 : _GEN_2766; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2896 = _T_6 ? mem_68 : _GEN_2767; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2897 = _T_6 ? mem_69 : _GEN_2768; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2898 = _T_6 ? mem_70 : _GEN_2769; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2899 = _T_6 ? mem_71 : _GEN_2770; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2900 = _T_6 ? mem_72 : _GEN_2771; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2901 = _T_6 ? mem_73 : _GEN_2772; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2902 = _T_6 ? mem_74 : _GEN_2773; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2903 = _T_6 ? mem_75 : _GEN_2774; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2904 = _T_6 ? mem_76 : _GEN_2775; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2905 = _T_6 ? mem_77 : _GEN_2776; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2906 = _T_6 ? mem_78 : _GEN_2777; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2907 = _T_6 ? mem_79 : _GEN_2778; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2908 = _T_6 ? mem_80 : _GEN_2779; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2909 = _T_6 ? mem_81 : _GEN_2780; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2910 = _T_6 ? mem_82 : _GEN_2781; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2911 = _T_6 ? mem_83 : _GEN_2782; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2912 = _T_6 ? mem_84 : _GEN_2783; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2913 = _T_6 ? mem_85 : _GEN_2784; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2914 = _T_6 ? mem_86 : _GEN_2785; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2915 = _T_6 ? mem_87 : _GEN_2786; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2916 = _T_6 ? mem_88 : _GEN_2787; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2917 = _T_6 ? mem_89 : _GEN_2788; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2918 = _T_6 ? mem_90 : _GEN_2789; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2919 = _T_6 ? mem_91 : _GEN_2790; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2920 = _T_6 ? mem_92 : _GEN_2791; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2921 = _T_6 ? mem_93 : _GEN_2792; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2922 = _T_6 ? mem_94 : _GEN_2793; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2923 = _T_6 ? mem_95 : _GEN_2794; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2924 = _T_6 ? mem_96 : _GEN_2795; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2925 = _T_6 ? mem_97 : _GEN_2796; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2926 = _T_6 ? mem_98 : _GEN_2797; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2927 = _T_6 ? mem_99 : _GEN_2798; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2928 = _T_6 ? mem_100 : _GEN_2799; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2929 = _T_6 ? mem_101 : _GEN_2800; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2930 = _T_6 ? mem_102 : _GEN_2801; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2931 = _T_6 ? mem_103 : _GEN_2802; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2932 = _T_6 ? mem_104 : _GEN_2803; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2933 = _T_6 ? mem_105 : _GEN_2804; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2934 = _T_6 ? mem_106 : _GEN_2805; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2935 = _T_6 ? mem_107 : _GEN_2806; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2936 = _T_6 ? mem_108 : _GEN_2807; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2937 = _T_6 ? mem_109 : _GEN_2808; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2938 = _T_6 ? mem_110 : _GEN_2809; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2939 = _T_6 ? mem_111 : _GEN_2810; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2940 = _T_6 ? mem_112 : _GEN_2811; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2941 = _T_6 ? mem_113 : _GEN_2812; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2942 = _T_6 ? mem_114 : _GEN_2813; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2943 = _T_6 ? mem_115 : _GEN_2814; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2944 = _T_6 ? mem_116 : _GEN_2815; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2945 = _T_6 ? mem_117 : _GEN_2816; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2946 = _T_6 ? mem_118 : _GEN_2817; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2947 = _T_6 ? mem_119 : _GEN_2818; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2948 = _T_6 ? mem_120 : _GEN_2819; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2949 = _T_6 ? mem_121 : _GEN_2820; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2950 = _T_6 ? mem_122 : _GEN_2821; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2951 = _T_6 ? mem_123 : _GEN_2822; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2952 = _T_6 ? mem_124 : _GEN_2823; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2953 = _T_6 ? mem_125 : _GEN_2824; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2954 = _T_6 ? mem_126 : _GEN_2825; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2955 = _T_6 ? mem_127 : _GEN_2826; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2956 = _T_5 ? 32'h0 : _GEN_2827; // @[Conditional.scala 39:67 data.scala 41:20]
  wire [31:0] _GEN_2957 = _T_5 ? mem_0 : _GEN_2828; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2958 = _T_5 ? mem_1 : _GEN_2829; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2959 = _T_5 ? mem_2 : _GEN_2830; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2960 = _T_5 ? mem_3 : _GEN_2831; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2961 = _T_5 ? mem_4 : _GEN_2832; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2962 = _T_5 ? mem_5 : _GEN_2833; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2963 = _T_5 ? mem_6 : _GEN_2834; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2964 = _T_5 ? mem_7 : _GEN_2835; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2965 = _T_5 ? mem_8 : _GEN_2836; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2966 = _T_5 ? mem_9 : _GEN_2837; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2967 = _T_5 ? mem_10 : _GEN_2838; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2968 = _T_5 ? mem_11 : _GEN_2839; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2969 = _T_5 ? mem_12 : _GEN_2840; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2970 = _T_5 ? mem_13 : _GEN_2841; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2971 = _T_5 ? mem_14 : _GEN_2842; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2972 = _T_5 ? mem_15 : _GEN_2843; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2973 = _T_5 ? mem_16 : _GEN_2844; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2974 = _T_5 ? mem_17 : _GEN_2845; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2975 = _T_5 ? mem_18 : _GEN_2846; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2976 = _T_5 ? mem_19 : _GEN_2847; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2977 = _T_5 ? mem_20 : _GEN_2848; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2978 = _T_5 ? mem_21 : _GEN_2849; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2979 = _T_5 ? mem_22 : _GEN_2850; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2980 = _T_5 ? mem_23 : _GEN_2851; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2981 = _T_5 ? mem_24 : _GEN_2852; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2982 = _T_5 ? mem_25 : _GEN_2853; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2983 = _T_5 ? mem_26 : _GEN_2854; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2984 = _T_5 ? mem_27 : _GEN_2855; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2985 = _T_5 ? mem_28 : _GEN_2856; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2986 = _T_5 ? mem_29 : _GEN_2857; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2987 = _T_5 ? mem_30 : _GEN_2858; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2988 = _T_5 ? mem_31 : _GEN_2859; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2989 = _T_5 ? mem_32 : _GEN_2860; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2990 = _T_5 ? mem_33 : _GEN_2861; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2991 = _T_5 ? mem_34 : _GEN_2862; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2992 = _T_5 ? mem_35 : _GEN_2863; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2993 = _T_5 ? mem_36 : _GEN_2864; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2994 = _T_5 ? mem_37 : _GEN_2865; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2995 = _T_5 ? mem_38 : _GEN_2866; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2996 = _T_5 ? mem_39 : _GEN_2867; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2997 = _T_5 ? mem_40 : _GEN_2868; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2998 = _T_5 ? mem_41 : _GEN_2869; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_2999 = _T_5 ? mem_42 : _GEN_2870; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3000 = _T_5 ? mem_43 : _GEN_2871; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3001 = _T_5 ? mem_44 : _GEN_2872; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3002 = _T_5 ? mem_45 : _GEN_2873; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3003 = _T_5 ? mem_46 : _GEN_2874; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3004 = _T_5 ? mem_47 : _GEN_2875; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3005 = _T_5 ? mem_48 : _GEN_2876; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3006 = _T_5 ? mem_49 : _GEN_2877; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3007 = _T_5 ? mem_50 : _GEN_2878; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3008 = _T_5 ? mem_51 : _GEN_2879; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3009 = _T_5 ? mem_52 : _GEN_2880; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3010 = _T_5 ? mem_53 : _GEN_2881; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3011 = _T_5 ? mem_54 : _GEN_2882; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3012 = _T_5 ? mem_55 : _GEN_2883; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3013 = _T_5 ? mem_56 : _GEN_2884; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3014 = _T_5 ? mem_57 : _GEN_2885; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3015 = _T_5 ? mem_58 : _GEN_2886; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3016 = _T_5 ? mem_59 : _GEN_2887; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3017 = _T_5 ? mem_60 : _GEN_2888; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3018 = _T_5 ? mem_61 : _GEN_2889; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3019 = _T_5 ? mem_62 : _GEN_2890; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3020 = _T_5 ? mem_63 : _GEN_2891; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3021 = _T_5 ? mem_64 : _GEN_2892; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3022 = _T_5 ? mem_65 : _GEN_2893; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3023 = _T_5 ? mem_66 : _GEN_2894; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3024 = _T_5 ? mem_67 : _GEN_2895; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3025 = _T_5 ? mem_68 : _GEN_2896; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3026 = _T_5 ? mem_69 : _GEN_2897; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3027 = _T_5 ? mem_70 : _GEN_2898; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3028 = _T_5 ? mem_71 : _GEN_2899; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3029 = _T_5 ? mem_72 : _GEN_2900; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3030 = _T_5 ? mem_73 : _GEN_2901; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3031 = _T_5 ? mem_74 : _GEN_2902; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3032 = _T_5 ? mem_75 : _GEN_2903; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3033 = _T_5 ? mem_76 : _GEN_2904; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3034 = _T_5 ? mem_77 : _GEN_2905; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3035 = _T_5 ? mem_78 : _GEN_2906; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3036 = _T_5 ? mem_79 : _GEN_2907; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3037 = _T_5 ? mem_80 : _GEN_2908; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3038 = _T_5 ? mem_81 : _GEN_2909; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3039 = _T_5 ? mem_82 : _GEN_2910; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3040 = _T_5 ? mem_83 : _GEN_2911; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3041 = _T_5 ? mem_84 : _GEN_2912; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3042 = _T_5 ? mem_85 : _GEN_2913; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3043 = _T_5 ? mem_86 : _GEN_2914; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3044 = _T_5 ? mem_87 : _GEN_2915; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3045 = _T_5 ? mem_88 : _GEN_2916; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3046 = _T_5 ? mem_89 : _GEN_2917; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3047 = _T_5 ? mem_90 : _GEN_2918; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3048 = _T_5 ? mem_91 : _GEN_2919; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3049 = _T_5 ? mem_92 : _GEN_2920; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3050 = _T_5 ? mem_93 : _GEN_2921; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3051 = _T_5 ? mem_94 : _GEN_2922; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3052 = _T_5 ? mem_95 : _GEN_2923; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3053 = _T_5 ? mem_96 : _GEN_2924; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3054 = _T_5 ? mem_97 : _GEN_2925; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3055 = _T_5 ? mem_98 : _GEN_2926; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3056 = _T_5 ? mem_99 : _GEN_2927; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3057 = _T_5 ? mem_100 : _GEN_2928; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3058 = _T_5 ? mem_101 : _GEN_2929; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3059 = _T_5 ? mem_102 : _GEN_2930; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3060 = _T_5 ? mem_103 : _GEN_2931; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3061 = _T_5 ? mem_104 : _GEN_2932; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3062 = _T_5 ? mem_105 : _GEN_2933; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3063 = _T_5 ? mem_106 : _GEN_2934; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3064 = _T_5 ? mem_107 : _GEN_2935; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3065 = _T_5 ? mem_108 : _GEN_2936; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3066 = _T_5 ? mem_109 : _GEN_2937; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3067 = _T_5 ? mem_110 : _GEN_2938; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3068 = _T_5 ? mem_111 : _GEN_2939; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3069 = _T_5 ? mem_112 : _GEN_2940; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3070 = _T_5 ? mem_113 : _GEN_2941; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3071 = _T_5 ? mem_114 : _GEN_2942; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3072 = _T_5 ? mem_115 : _GEN_2943; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3073 = _T_5 ? mem_116 : _GEN_2944; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3074 = _T_5 ? mem_117 : _GEN_2945; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3075 = _T_5 ? mem_118 : _GEN_2946; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3076 = _T_5 ? mem_119 : _GEN_2947; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3077 = _T_5 ? mem_120 : _GEN_2948; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3078 = _T_5 ? mem_121 : _GEN_2949; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3079 = _T_5 ? mem_122 : _GEN_2950; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3080 = _T_5 ? mem_123 : _GEN_2951; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3081 = _T_5 ? mem_124 : _GEN_2952; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3082 = _T_5 ? mem_125 : _GEN_2953; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3083 = _T_5 ? mem_126 : _GEN_2954; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3084 = _T_5 ? mem_127 : _GEN_2955; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3085 = _T_4 ? 32'h0 : _GEN_2956; // @[Conditional.scala 39:67 data.scala 38:20]
  wire [31:0] _GEN_3086 = _T_4 ? mem_0 : _GEN_2957; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3087 = _T_4 ? mem_1 : _GEN_2958; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3088 = _T_4 ? mem_2 : _GEN_2959; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3089 = _T_4 ? mem_3 : _GEN_2960; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3090 = _T_4 ? mem_4 : _GEN_2961; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3091 = _T_4 ? mem_5 : _GEN_2962; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3092 = _T_4 ? mem_6 : _GEN_2963; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3093 = _T_4 ? mem_7 : _GEN_2964; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3094 = _T_4 ? mem_8 : _GEN_2965; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3095 = _T_4 ? mem_9 : _GEN_2966; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3096 = _T_4 ? mem_10 : _GEN_2967; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3097 = _T_4 ? mem_11 : _GEN_2968; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3098 = _T_4 ? mem_12 : _GEN_2969; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3099 = _T_4 ? mem_13 : _GEN_2970; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3100 = _T_4 ? mem_14 : _GEN_2971; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3101 = _T_4 ? mem_15 : _GEN_2972; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3102 = _T_4 ? mem_16 : _GEN_2973; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3103 = _T_4 ? mem_17 : _GEN_2974; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3104 = _T_4 ? mem_18 : _GEN_2975; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3105 = _T_4 ? mem_19 : _GEN_2976; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3106 = _T_4 ? mem_20 : _GEN_2977; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3107 = _T_4 ? mem_21 : _GEN_2978; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3108 = _T_4 ? mem_22 : _GEN_2979; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3109 = _T_4 ? mem_23 : _GEN_2980; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3110 = _T_4 ? mem_24 : _GEN_2981; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3111 = _T_4 ? mem_25 : _GEN_2982; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3112 = _T_4 ? mem_26 : _GEN_2983; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3113 = _T_4 ? mem_27 : _GEN_2984; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3114 = _T_4 ? mem_28 : _GEN_2985; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3115 = _T_4 ? mem_29 : _GEN_2986; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3116 = _T_4 ? mem_30 : _GEN_2987; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3117 = _T_4 ? mem_31 : _GEN_2988; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3118 = _T_4 ? mem_32 : _GEN_2989; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3119 = _T_4 ? mem_33 : _GEN_2990; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3120 = _T_4 ? mem_34 : _GEN_2991; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3121 = _T_4 ? mem_35 : _GEN_2992; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3122 = _T_4 ? mem_36 : _GEN_2993; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3123 = _T_4 ? mem_37 : _GEN_2994; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3124 = _T_4 ? mem_38 : _GEN_2995; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3125 = _T_4 ? mem_39 : _GEN_2996; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3126 = _T_4 ? mem_40 : _GEN_2997; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3127 = _T_4 ? mem_41 : _GEN_2998; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3128 = _T_4 ? mem_42 : _GEN_2999; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3129 = _T_4 ? mem_43 : _GEN_3000; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3130 = _T_4 ? mem_44 : _GEN_3001; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3131 = _T_4 ? mem_45 : _GEN_3002; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3132 = _T_4 ? mem_46 : _GEN_3003; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3133 = _T_4 ? mem_47 : _GEN_3004; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3134 = _T_4 ? mem_48 : _GEN_3005; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3135 = _T_4 ? mem_49 : _GEN_3006; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3136 = _T_4 ? mem_50 : _GEN_3007; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3137 = _T_4 ? mem_51 : _GEN_3008; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3138 = _T_4 ? mem_52 : _GEN_3009; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3139 = _T_4 ? mem_53 : _GEN_3010; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3140 = _T_4 ? mem_54 : _GEN_3011; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3141 = _T_4 ? mem_55 : _GEN_3012; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3142 = _T_4 ? mem_56 : _GEN_3013; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3143 = _T_4 ? mem_57 : _GEN_3014; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3144 = _T_4 ? mem_58 : _GEN_3015; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3145 = _T_4 ? mem_59 : _GEN_3016; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3146 = _T_4 ? mem_60 : _GEN_3017; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3147 = _T_4 ? mem_61 : _GEN_3018; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3148 = _T_4 ? mem_62 : _GEN_3019; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3149 = _T_4 ? mem_63 : _GEN_3020; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3150 = _T_4 ? mem_64 : _GEN_3021; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3151 = _T_4 ? mem_65 : _GEN_3022; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3152 = _T_4 ? mem_66 : _GEN_3023; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3153 = _T_4 ? mem_67 : _GEN_3024; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3154 = _T_4 ? mem_68 : _GEN_3025; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3155 = _T_4 ? mem_69 : _GEN_3026; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3156 = _T_4 ? mem_70 : _GEN_3027; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3157 = _T_4 ? mem_71 : _GEN_3028; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3158 = _T_4 ? mem_72 : _GEN_3029; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3159 = _T_4 ? mem_73 : _GEN_3030; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3160 = _T_4 ? mem_74 : _GEN_3031; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3161 = _T_4 ? mem_75 : _GEN_3032; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3162 = _T_4 ? mem_76 : _GEN_3033; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3163 = _T_4 ? mem_77 : _GEN_3034; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3164 = _T_4 ? mem_78 : _GEN_3035; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3165 = _T_4 ? mem_79 : _GEN_3036; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3166 = _T_4 ? mem_80 : _GEN_3037; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3167 = _T_4 ? mem_81 : _GEN_3038; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3168 = _T_4 ? mem_82 : _GEN_3039; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3169 = _T_4 ? mem_83 : _GEN_3040; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3170 = _T_4 ? mem_84 : _GEN_3041; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3171 = _T_4 ? mem_85 : _GEN_3042; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3172 = _T_4 ? mem_86 : _GEN_3043; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3173 = _T_4 ? mem_87 : _GEN_3044; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3174 = _T_4 ? mem_88 : _GEN_3045; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3175 = _T_4 ? mem_89 : _GEN_3046; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3176 = _T_4 ? mem_90 : _GEN_3047; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3177 = _T_4 ? mem_91 : _GEN_3048; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3178 = _T_4 ? mem_92 : _GEN_3049; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3179 = _T_4 ? mem_93 : _GEN_3050; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3180 = _T_4 ? mem_94 : _GEN_3051; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3181 = _T_4 ? mem_95 : _GEN_3052; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3182 = _T_4 ? mem_96 : _GEN_3053; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3183 = _T_4 ? mem_97 : _GEN_3054; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3184 = _T_4 ? mem_98 : _GEN_3055; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3185 = _T_4 ? mem_99 : _GEN_3056; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3186 = _T_4 ? mem_100 : _GEN_3057; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3187 = _T_4 ? mem_101 : _GEN_3058; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3188 = _T_4 ? mem_102 : _GEN_3059; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3189 = _T_4 ? mem_103 : _GEN_3060; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3190 = _T_4 ? mem_104 : _GEN_3061; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3191 = _T_4 ? mem_105 : _GEN_3062; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3192 = _T_4 ? mem_106 : _GEN_3063; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3193 = _T_4 ? mem_107 : _GEN_3064; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3194 = _T_4 ? mem_108 : _GEN_3065; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3195 = _T_4 ? mem_109 : _GEN_3066; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3196 = _T_4 ? mem_110 : _GEN_3067; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3197 = _T_4 ? mem_111 : _GEN_3068; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3198 = _T_4 ? mem_112 : _GEN_3069; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3199 = _T_4 ? mem_113 : _GEN_3070; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3200 = _T_4 ? mem_114 : _GEN_3071; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3201 = _T_4 ? mem_115 : _GEN_3072; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3202 = _T_4 ? mem_116 : _GEN_3073; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3203 = _T_4 ? mem_117 : _GEN_3074; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3204 = _T_4 ? mem_118 : _GEN_3075; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3205 = _T_4 ? mem_119 : _GEN_3076; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3206 = _T_4 ? mem_120 : _GEN_3077; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3207 = _T_4 ? mem_121 : _GEN_3078; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3208 = _T_4 ? mem_122 : _GEN_3079; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3209 = _T_4 ? mem_123 : _GEN_3080; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3210 = _T_4 ? mem_124 : _GEN_3081; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3211 = _T_4 ? mem_125 : _GEN_3082; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3212 = _T_4 ? mem_126 : _GEN_3083; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3213 = _T_4 ? mem_127 : _GEN_3084; // @[Conditional.scala 39:67 data.scala 18:16]
  wire [31:0] _GEN_3214 = _T_3 ? 32'h0 : _GEN_3085; // @[Conditional.scala 39:67 data.scala 35:20]
  wire [31:0] _GEN_3343 = _T_2 ? 32'h0 : _GEN_3214; // @[Conditional.scala 39:67 data.scala 32:20]
  wire [31:0] _GEN_3472 = _T_1 ? 32'h0 : _GEN_3343; // @[Conditional.scala 40:58 data.scala 29:20]
  assign io_data_read = reset ? 32'h0 : _GEN_3472; // @[data.scala 21:3 data.scala 16:16]
  always @(posedge clock) begin
    if (reset) begin // @[data.scala 21:3]
      mem_0 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_0 <= _GEN_3086;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_1 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_1 <= _GEN_3087;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_2 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_2 <= _GEN_3088;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_3 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_3 <= _GEN_3089;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_4 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_4 <= _GEN_3090;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_5 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_5 <= _GEN_3091;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_6 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_6 <= _GEN_3092;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_7 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_7 <= _GEN_3093;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_8 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_8 <= _GEN_3094;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_9 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_9 <= _GEN_3095;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_10 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_10 <= _GEN_3096;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_11 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_11 <= _GEN_3097;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_12 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_12 <= _GEN_3098;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_13 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_13 <= _GEN_3099;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_14 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_14 <= _GEN_3100;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_15 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_15 <= _GEN_3101;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_16 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_16 <= _GEN_3102;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_17 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_17 <= _GEN_3103;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_18 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_18 <= _GEN_3104;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_19 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_19 <= _GEN_3105;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_20 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_20 <= _GEN_3106;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_21 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_21 <= _GEN_3107;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_22 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_22 <= _GEN_3108;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_23 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_23 <= _GEN_3109;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_24 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_24 <= _GEN_3110;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_25 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_25 <= _GEN_3111;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_26 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_26 <= _GEN_3112;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_27 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_27 <= _GEN_3113;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_28 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_28 <= _GEN_3114;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_29 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_29 <= _GEN_3115;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_30 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_30 <= _GEN_3116;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_31 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_31 <= _GEN_3117;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_32 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_32 <= _GEN_3118;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_33 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_33 <= _GEN_3119;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_34 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_34 <= _GEN_3120;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_35 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_35 <= _GEN_3121;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_36 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_36 <= _GEN_3122;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_37 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_37 <= _GEN_3123;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_38 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_38 <= _GEN_3124;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_39 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_39 <= _GEN_3125;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_40 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_40 <= _GEN_3126;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_41 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_41 <= _GEN_3127;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_42 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_42 <= _GEN_3128;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_43 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_43 <= _GEN_3129;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_44 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_44 <= _GEN_3130;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_45 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_45 <= _GEN_3131;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_46 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_46 <= _GEN_3132;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_47 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_47 <= _GEN_3133;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_48 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_48 <= _GEN_3134;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_49 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_49 <= _GEN_3135;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_50 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_50 <= _GEN_3136;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_51 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_51 <= _GEN_3137;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_52 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_52 <= _GEN_3138;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_53 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_53 <= _GEN_3139;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_54 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_54 <= _GEN_3140;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_55 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_55 <= _GEN_3141;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_56 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_56 <= _GEN_3142;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_57 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_57 <= _GEN_3143;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_58 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_58 <= _GEN_3144;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_59 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_59 <= _GEN_3145;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_60 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_60 <= _GEN_3146;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_61 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_61 <= _GEN_3147;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_62 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_62 <= _GEN_3148;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_63 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_63 <= _GEN_3149;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_64 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_64 <= _GEN_3150;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_65 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_65 <= _GEN_3151;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_66 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_66 <= _GEN_3152;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_67 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_67 <= _GEN_3153;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_68 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_68 <= _GEN_3154;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_69 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_69 <= _GEN_3155;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_70 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_70 <= _GEN_3156;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_71 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_71 <= _GEN_3157;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_72 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_72 <= _GEN_3158;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_73 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_73 <= _GEN_3159;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_74 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_74 <= _GEN_3160;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_75 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_75 <= _GEN_3161;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_76 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_76 <= _GEN_3162;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_77 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_77 <= _GEN_3163;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_78 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_78 <= _GEN_3164;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_79 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_79 <= _GEN_3165;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_80 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_80 <= _GEN_3166;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_81 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_81 <= _GEN_3167;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_82 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_82 <= _GEN_3168;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_83 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_83 <= _GEN_3169;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_84 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_84 <= _GEN_3170;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_85 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_85 <= _GEN_3171;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_86 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_86 <= _GEN_3172;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_87 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_87 <= _GEN_3173;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_88 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_88 <= _GEN_3174;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_89 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_89 <= _GEN_3175;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_90 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_90 <= _GEN_3176;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_91 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_91 <= _GEN_3177;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_92 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_92 <= _GEN_3178;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_93 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_93 <= _GEN_3179;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_94 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_94 <= _GEN_3180;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_95 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_95 <= _GEN_3181;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_96 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_96 <= _GEN_3182;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_97 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_97 <= _GEN_3183;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_98 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_98 <= _GEN_3184;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_99 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_99 <= _GEN_3185;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_100 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_100 <= _GEN_3186;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_101 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_101 <= _GEN_3187;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_102 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_102 <= _GEN_3188;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_103 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_103 <= _GEN_3189;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_104 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_104 <= _GEN_3190;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_105 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_105 <= _GEN_3191;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_106 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_106 <= _GEN_3192;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_107 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_107 <= _GEN_3193;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_108 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_108 <= _GEN_3194;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_109 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_109 <= _GEN_3195;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_110 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_110 <= _GEN_3196;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_111 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_111 <= _GEN_3197;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_112 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_112 <= _GEN_3198;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_113 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_113 <= _GEN_3199;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_114 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_114 <= _GEN_3200;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_115 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_115 <= _GEN_3201;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_116 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_116 <= _GEN_3202;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_117 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_117 <= _GEN_3203;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_118 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_118 <= _GEN_3204;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_119 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_119 <= _GEN_3205;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_120 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_120 <= _GEN_3206;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_121 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_121 <= _GEN_3207;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_122 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_122 <= _GEN_3208;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_123 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_123 <= _GEN_3209;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_124 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_124 <= _GEN_3210;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_125 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_125 <= _GEN_3211;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_126 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_126 <= _GEN_3212;
        end
      end
    end
    if (reset) begin // @[data.scala 21:3]
      mem_127 <= 32'h0; // @[data.scala 23:14]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          mem_127 <= _GEN_3213;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mem_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mem_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mem_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mem_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mem_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mem_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mem_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mem_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  mem_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mem_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mem_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mem_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mem_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mem_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mem_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mem_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  mem_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  mem_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  mem_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mem_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mem_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mem_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mem_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mem_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mem_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mem_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mem_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mem_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mem_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mem_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mem_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mem_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mem_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mem_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mem_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mem_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mem_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mem_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mem_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mem_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mem_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mem_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mem_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mem_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mem_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mem_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mem_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mem_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mem_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mem_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mem_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mem_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mem_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mem_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mem_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mem_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mem_64 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mem_65 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mem_66 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mem_67 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mem_68 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mem_69 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mem_70 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mem_71 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mem_72 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mem_73 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mem_74 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mem_75 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mem_76 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mem_77 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mem_78 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mem_79 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mem_80 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mem_81 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mem_82 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mem_83 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mem_84 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mem_85 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mem_86 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mem_87 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mem_88 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mem_89 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mem_90 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mem_91 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mem_92 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mem_93 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mem_94 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mem_95 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mem_96 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mem_97 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mem_98 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mem_99 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mem_100 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mem_101 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mem_102 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mem_103 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mem_104 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mem_105 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mem_106 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mem_107 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mem_108 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mem_109 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mem_110 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mem_111 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mem_112 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mem_113 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mem_114 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mem_115 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mem_116 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mem_117 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mem_118 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mem_119 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mem_120 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mem_121 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mem_122 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mem_123 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mem_124 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mem_125 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mem_126 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mem_127 = _RAND_127[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module imm_gen(
  input  [7:0]  io_imm_ctrl,
  input  [31:0] io_instruction,
  output [31:0] io_imm
);
  wire  _T = 8'h8 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_14 = {io_instruction[31:12], 12'h0}; // @[imm_gen.scala 19:39]
  wire [34:0] _io_imm_T_1 = {{3'd0}, _GEN_14}; // @[imm_gen.scala 19:39]
  wire  _T_1 = 8'h1 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire  _T_3 = ~io_instruction[31]; // @[imm_gen.scala 22:31]
  wire [11:0] _GEN_15 = {io_instruction[7], 11'h0}; // @[imm_gen.scala 23:37]
  wire [15:0] _io_imm_T_3 = {{4'd0}, _GEN_15}; // @[imm_gen.scala 23:37]
  wire [10:0] _GEN_16 = {io_instruction[30:25], 5'h0}; // @[imm_gen.scala 23:69]
  wire [12:0] _io_imm_T_5 = {{2'd0}, _GEN_16}; // @[imm_gen.scala 23:69]
  wire [15:0] _GEN_17 = {{3'd0}, _io_imm_T_5}; // @[imm_gen.scala 23:45]
  wire [15:0] _io_imm_T_7 = _io_imm_T_3 + _GEN_17; // @[imm_gen.scala 23:45]
  wire [4:0] _io_imm_T_9 = {io_instruction[11:8], 1'h0}; // @[imm_gen.scala 23:99]
  wire [15:0] _GEN_18 = {{11'd0}, _io_imm_T_9}; // @[imm_gen.scala 23:76]
  wire [15:0] _io_imm_T_11 = _io_imm_T_7 + _GEN_18; // @[imm_gen.scala 23:76]
  wire [31:0] _GEN_23 = {{16'd0}, _io_imm_T_11}; // @[imm_gen.scala 26:106]
  wire [31:0] _io_imm_T_23 = _GEN_23 + 32'hffffffff; // @[imm_gen.scala 26:106]
  wire [43:0] _GEN_24 = {_io_imm_T_23, 12'h0}; // @[imm_gen.scala 26:121]
  wire [46:0] _io_imm_T_24 = {{3'd0}, _GEN_24}; // @[imm_gen.scala 26:121]
  wire [46:0] _GEN_0 = ~io_instruction[31] ? {{31'd0}, _io_imm_T_11} : _io_imm_T_24; // @[imm_gen.scala 22:39 imm_gen.scala 23:16 imm_gen.scala 26:16]
  wire  _T_4 = 8'h2 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire  _T_5 = 8'h0 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire  _T_6 = 8'h5 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire [19:0] _GEN_25 = {io_instruction[19:12], 12'h0}; // @[imm_gen.scala 37:41]
  wire [22:0] _io_imm_T_28 = {{3'd0}, _GEN_25}; // @[imm_gen.scala 37:41]
  wire [11:0] _GEN_26 = {io_instruction[20], 11'h0}; // @[imm_gen.scala 37:70]
  wire [15:0] _io_imm_T_30 = {{4'd0}, _GEN_26}; // @[imm_gen.scala 37:70]
  wire [22:0] _GEN_27 = {{7'd0}, _io_imm_T_30}; // @[imm_gen.scala 37:49]
  wire [22:0] _io_imm_T_32 = _io_imm_T_28 + _GEN_27; // @[imm_gen.scala 37:49]
  wire [10:0] _io_imm_T_34 = {io_instruction[30:21], 1'h0}; // @[imm_gen.scala 37:102]
  wire [22:0] _GEN_28 = {{12'd0}, _io_imm_T_34}; // @[imm_gen.scala 37:78]
  wire [22:0] _io_imm_T_36 = _io_imm_T_32 + _GEN_28; // @[imm_gen.scala 37:78]
  wire [31:0] _GEN_33 = {{9'd0}, _io_imm_T_36}; // @[imm_gen.scala 39:109]
  wire [31:0] _io_imm_T_48 = _GEN_33 + 32'hffffffff; // @[imm_gen.scala 39:109]
  wire [43:0] _GEN_34 = {_io_imm_T_48, 12'h0}; // @[imm_gen.scala 39:124]
  wire [46:0] _io_imm_T_49 = {{3'd0}, _GEN_34}; // @[imm_gen.scala 39:124]
  wire [46:0] _GEN_1 = _T_3 ? {{24'd0}, _io_imm_T_36} : _io_imm_T_49; // @[imm_gen.scala 36:39 imm_gen.scala 37:16 imm_gen.scala 39:16]
  wire  _T_9 = 8'h3 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire [46:0] _GEN_35 = {{35'd0}, io_instruction[31:20]}; // @[imm_gen.scala 47:41]
  wire [46:0] _io_imm_T_54 = _GEN_35 + 47'h7fffffff800; // @[imm_gen.scala 47:41]
  wire [46:0] _GEN_2 = _T_3 ? {{35'd0}, io_instruction[31:20]} : _io_imm_T_54; // @[imm_gen.scala 43:39 imm_gen.scala 44:16 imm_gen.scala 47:16]
  wire  _T_12 = 8'h4 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire  _T_15 = 8'h9 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire  _T_16 = 8'h6 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire  _T_17 = 8'h7 == io_imm_ctrl; // @[Conditional.scala 37:30]
  wire [11:0] _GEN_38 = {io_instruction[31:25], 5'h0}; // @[imm_gen.scala 65:39]
  wire [13:0] _io_imm_T_63 = {{2'd0}, _GEN_38}; // @[imm_gen.scala 65:39]
  wire [13:0] _GEN_39 = {{9'd0}, io_instruction[11:7]}; // @[imm_gen.scala 65:46]
  wire [13:0] _io_imm_T_66 = _io_imm_T_63 + _GEN_39; // @[imm_gen.scala 65:46]
  wire [13:0] _GEN_4 = _T_17 ? _io_imm_T_66 : 14'h0; // @[Conditional.scala 39:67 imm_gen.scala 65:14 imm_gen.scala 15:10]
  wire [13:0] _GEN_5 = _T_16 ? 14'h0 : _GEN_4; // @[Conditional.scala 39:67 imm_gen.scala 62:14]
  wire [34:0] _GEN_6 = _T_15 ? _io_imm_T_1 : {{21'd0}, _GEN_5}; // @[Conditional.scala 39:67 imm_gen.scala 59:14]
  wire [46:0] _GEN_7 = _T_12 ? _GEN_2 : {{12'd0}, _GEN_6}; // @[Conditional.scala 39:67]
  wire [46:0] _GEN_8 = _T_9 ? _GEN_2 : _GEN_7; // @[Conditional.scala 39:67]
  wire [46:0] _GEN_9 = _T_6 ? _GEN_1 : _GEN_8; // @[Conditional.scala 39:67]
  wire [46:0] _GEN_10 = _T_5 ? {{35'd0}, io_instruction[31:20]} : _GEN_9; // @[Conditional.scala 39:67 imm_gen.scala 33:14]
  wire [46:0] _GEN_11 = _T_4 ? {{42'd0}, io_instruction[24:20]} : _GEN_10; // @[Conditional.scala 39:67 imm_gen.scala 30:14]
  wire [46:0] _GEN_12 = _T_1 ? _GEN_0 : _GEN_11; // @[Conditional.scala 39:67]
  wire [46:0] _GEN_13 = _T ? {{12'd0}, _io_imm_T_1} : _GEN_12; // @[Conditional.scala 40:58 imm_gen.scala 19:14]
  assign io_imm = _GEN_13[31:0];
endmodule
module instruction(
  input         reset,
  input  [31:0] io_pc,
  output [31:0] io_instruction
);
  wire [31:0] _io_instruction_T = io_pc / 3'h4; // @[instruction.scala 98:36]
  wire [31:0] _GEN_1 = 7'h1 == _io_instruction_T[6:0] ? 32'h3fb95ab7 : 32'h18f06a13; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_2 = 7'h2 == _io_instruction_T[6:0] ? 32'h15a6a33 : _GEN_1; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_3 = 7'h3 == _io_instruction_T[6:0] ? 32'h98765ab7 : _GEN_2; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_4 = 7'h4 == _io_instruction_T[6:0] ? 32'h345a8a93 : _GEN_3; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_5 = 7'h5 == _io_instruction_T[6:0] ? 32'hc00a0b13 : _GEN_4; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_6 = 7'h6 == _io_instruction_T[6:0] ? 32'h7bca4b93 : _GEN_5; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_7 = 7'h7 == _io_instruction_T[6:0] ? 32'h34a3b13 : _GEN_6; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_8 = 7'h8 == _io_instruction_T[6:0] ? 32'hfffa3b93 : _GEN_7; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_9 = 7'h9 == _io_instruction_T[6:0] ? 32'h765a7b13 : _GEN_8; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_10 = 7'ha == _io_instruction_T[6:0] ? 32'hfffa2b93 : _GEN_9; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_11 = 7'hb == _io_instruction_T[6:0] ? 32'h414a8b33 : _GEN_10; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_12 = 7'hc == _io_instruction_T[6:0] ? 32'h16a4bb3 : _GEN_11; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_13 = 7'hd == _io_instruction_T[6:0] ? 32'h14a8b33 : _GEN_12; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_14 = 7'he == _io_instruction_T[6:0] ? 32'h414b0b33 : _GEN_13; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_15 = 7'hf == _io_instruction_T[6:0] ? 32'h16bebb3 : _GEN_14; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_16 = 7'h10 == _io_instruction_T[6:0] ? 32'h16bfbb3 : _GEN_15; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_17 = 7'h11 == _io_instruction_T[6:0] ? 32'h15a2b33 : _GEN_16; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_18 = 7'h12 == _io_instruction_T[6:0] ? 32'h15a3bb3 : _GEN_17; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_19 = 7'h13 == _io_instruction_T[6:0] ? 32'h418193 : _GEN_18; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_20 = 7'h14 == _io_instruction_T[6:0] ? 32'h3a1b33 : _GEN_19; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_21 = 7'h15 == _io_instruction_T[6:0] ? 32'h3adb33 : _GEN_20; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_22 = 7'h16 == _io_instruction_T[6:0] ? 32'h403adb33 : _GEN_21; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_23 = 7'h17 == _io_instruction_T[6:0] ? 32'h10a9b93 : _GEN_22; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_24 = 7'h18 == _io_instruction_T[6:0] ? 32'h8adb93 : _GEN_23; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_25 = 7'h19 == _io_instruction_T[6:0] ? 32'h408adb93 : _GEN_24; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_26 = 7'h1a == _io_instruction_T[6:0] ? 32'h193 : _GEN_25; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_27 = 7'h1b == _io_instruction_T[6:0] ? 32'hf500293 : _GEN_26; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_28 = 7'h1c == _io_instruction_T[6:0] ? 32'h141a023 : _GEN_27; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_29 = 7'h1d == _io_instruction_T[6:0] ? 32'h151a223 : _GEN_28; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_30 = 7'h1e == _io_instruction_T[6:0] ? 32'h171a423 : _GEN_29; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_31 = 7'h1f == _io_instruction_T[6:0] ? 32'h1619223 : _GEN_30; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_32 = 7'h20 == _io_instruction_T[6:0] ? 32'h1419523 : _GEN_31; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_33 = 7'h21 == _io_instruction_T[6:0] ? 32'h5183a3 : _GEN_32; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_34 = 7'h22 == _io_instruction_T[6:0] ? 32'h5184a3 : _GEN_33; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_35 = 7'h23 == _io_instruction_T[6:0] ? 32'h518423 : _GEN_34; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_36 = 7'h24 == _io_instruction_T[6:0] ? 32'h1ab03 : _GEN_35; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_37 = 7'h25 == _io_instruction_T[6:0] ? 32'h161a623 : _GEN_36; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_38 = 7'h26 == _io_instruction_T[6:0] ? 32'h819b83 : _GEN_37; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_39 = 7'h27 == _io_instruction_T[6:0] ? 32'h171a823 : _GEN_38; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_40 = 7'h28 == _io_instruction_T[6:0] ? 32'h81db83 : _GEN_39; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_41 = 7'h29 == _io_instruction_T[6:0] ? 32'h141aa23 : _GEN_40; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_42 = 7'h2a == _io_instruction_T[6:0] ? 32'h718b03 : _GEN_41; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_43 = 7'h2b == _io_instruction_T[6:0] ? 32'h151ac23 : _GEN_42; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_44 = 7'h2c == _io_instruction_T[6:0] ? 32'h71cb83 : _GEN_43; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_45 = 7'h2d == _io_instruction_T[6:0] ? 32'h171ae23 : _GEN_44; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_46 = 7'h2e == _io_instruction_T[6:0] ? 32'h181cb83 : _GEN_45; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_47 = 7'h2f == _io_instruction_T[6:0] ? 32'h371a023 : _GEN_46; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_48 = 7'h30 == _io_instruction_T[6:0] ? 32'h1a223 : _GEN_47; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_49 = 7'h31 == _io_instruction_T[6:0] ? 32'h9074b3 : _GEN_48; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_50 = 7'h32 == _io_instruction_T[6:0] ? 32'h15a1463 : _GEN_49; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_51 = 7'h33 == _io_instruction_T[6:0] ? 32'h148493 : _GEN_50; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_52 = 7'h34 == _io_instruction_T[6:0] ? 32'h15a5463 : _GEN_51; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_53 = 7'h35 == _io_instruction_T[6:0] ? 32'h148493 : _GEN_52; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_54 = 7'h36 == _io_instruction_T[6:0] ? 32'h15a7463 : _GEN_53; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_55 = 7'h37 == _io_instruction_T[6:0] ? 32'h248493 : _GEN_54; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_56 = 7'h38 == _io_instruction_T[6:0] ? 32'h15a4463 : _GEN_55; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_57 = 7'h39 == _io_instruction_T[6:0] ? 32'h348493 : _GEN_56; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_58 = 7'h3a == _io_instruction_T[6:0] ? 32'h15a6463 : _GEN_57; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_59 = 7'h3b == _io_instruction_T[6:0] ? 32'h448493 : _GEN_58; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_60 = 7'h3c == _io_instruction_T[6:0] ? 32'h181ac83 : _GEN_59; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_61 = 7'h3d == _io_instruction_T[6:0] ? 32'h19a8463 : _GEN_60; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_62 = 7'h3e == _io_instruction_T[6:0] ? 32'h548493 : _GEN_61; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_63 = 7'h3f == _io_instruction_T[6:0] ? 32'h91a223 : _GEN_62; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_64 = 7'h40 == _io_instruction_T[6:0] ? 32'h41a503 : _GEN_63; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_65 = 7'h41 == _io_instruction_T[6:0] ? 32'hc000ef : _GEN_64; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_66 = 7'h42 == _io_instruction_T[6:0] ? 32'h850513 : _GEN_65; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_67 = 7'h43 == _io_instruction_T[6:0] ? 32'ha1a223 : _GEN_66; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_68 = 7'h44 == _io_instruction_T[6:0] ? 32'h45c56513 : _GEN_67; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_69 = 7'h45 == _io_instruction_T[6:0] ? 32'ha1a223 : _GEN_68; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_70 = 7'h46 == _io_instruction_T[6:0] ? 32'h8067 : _GEN_69; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_71 = 7'h47 == _io_instruction_T[6:0] ? 32'h0 : _GEN_70; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_72 = 7'h48 == _io_instruction_T[6:0] ? 32'h0 : _GEN_71; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_73 = 7'h49 == _io_instruction_T[6:0] ? 32'h0 : _GEN_72; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_74 = 7'h4a == _io_instruction_T[6:0] ? 32'h0 : _GEN_73; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_75 = 7'h4b == _io_instruction_T[6:0] ? 32'h0 : _GEN_74; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_76 = 7'h4c == _io_instruction_T[6:0] ? 32'h0 : _GEN_75; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_77 = 7'h4d == _io_instruction_T[6:0] ? 32'h0 : _GEN_76; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_78 = 7'h4e == _io_instruction_T[6:0] ? 32'h0 : _GEN_77; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_79 = 7'h4f == _io_instruction_T[6:0] ? 32'h0 : _GEN_78; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_80 = 7'h50 == _io_instruction_T[6:0] ? 32'h0 : _GEN_79; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_81 = 7'h51 == _io_instruction_T[6:0] ? 32'h0 : _GEN_80; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_82 = 7'h52 == _io_instruction_T[6:0] ? 32'h0 : _GEN_81; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_83 = 7'h53 == _io_instruction_T[6:0] ? 32'h0 : _GEN_82; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_84 = 7'h54 == _io_instruction_T[6:0] ? 32'h0 : _GEN_83; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_85 = 7'h55 == _io_instruction_T[6:0] ? 32'h0 : _GEN_84; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_86 = 7'h56 == _io_instruction_T[6:0] ? 32'h0 : _GEN_85; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_87 = 7'h57 == _io_instruction_T[6:0] ? 32'h0 : _GEN_86; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_88 = 7'h58 == _io_instruction_T[6:0] ? 32'h0 : _GEN_87; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_89 = 7'h59 == _io_instruction_T[6:0] ? 32'h0 : _GEN_88; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_90 = 7'h5a == _io_instruction_T[6:0] ? 32'h0 : _GEN_89; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_91 = 7'h5b == _io_instruction_T[6:0] ? 32'h0 : _GEN_90; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_92 = 7'h5c == _io_instruction_T[6:0] ? 32'h0 : _GEN_91; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_93 = 7'h5d == _io_instruction_T[6:0] ? 32'h0 : _GEN_92; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_94 = 7'h5e == _io_instruction_T[6:0] ? 32'h0 : _GEN_93; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_95 = 7'h5f == _io_instruction_T[6:0] ? 32'h0 : _GEN_94; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_96 = 7'h60 == _io_instruction_T[6:0] ? 32'h0 : _GEN_95; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_97 = 7'h61 == _io_instruction_T[6:0] ? 32'h0 : _GEN_96; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_98 = 7'h62 == _io_instruction_T[6:0] ? 32'h0 : _GEN_97; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_99 = 7'h63 == _io_instruction_T[6:0] ? 32'h0 : _GEN_98; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_100 = 7'h64 == _io_instruction_T[6:0] ? 32'h0 : _GEN_99; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_101 = 7'h65 == _io_instruction_T[6:0] ? 32'h0 : _GEN_100; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_102 = 7'h66 == _io_instruction_T[6:0] ? 32'h0 : _GEN_101; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_103 = 7'h67 == _io_instruction_T[6:0] ? 32'h0 : _GEN_102; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_104 = 7'h68 == _io_instruction_T[6:0] ? 32'h0 : _GEN_103; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_105 = 7'h69 == _io_instruction_T[6:0] ? 32'h0 : _GEN_104; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_106 = 7'h6a == _io_instruction_T[6:0] ? 32'h0 : _GEN_105; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_107 = 7'h6b == _io_instruction_T[6:0] ? 32'h0 : _GEN_106; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_108 = 7'h6c == _io_instruction_T[6:0] ? 32'h0 : _GEN_107; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_109 = 7'h6d == _io_instruction_T[6:0] ? 32'h0 : _GEN_108; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_110 = 7'h6e == _io_instruction_T[6:0] ? 32'h0 : _GEN_109; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_111 = 7'h6f == _io_instruction_T[6:0] ? 32'h0 : _GEN_110; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_112 = 7'h70 == _io_instruction_T[6:0] ? 32'h0 : _GEN_111; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_113 = 7'h71 == _io_instruction_T[6:0] ? 32'h0 : _GEN_112; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_114 = 7'h72 == _io_instruction_T[6:0] ? 32'h0 : _GEN_113; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_115 = 7'h73 == _io_instruction_T[6:0] ? 32'h0 : _GEN_114; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_116 = 7'h74 == _io_instruction_T[6:0] ? 32'h0 : _GEN_115; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_117 = 7'h75 == _io_instruction_T[6:0] ? 32'h0 : _GEN_116; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_118 = 7'h76 == _io_instruction_T[6:0] ? 32'h0 : _GEN_117; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_119 = 7'h77 == _io_instruction_T[6:0] ? 32'h0 : _GEN_118; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_120 = 7'h78 == _io_instruction_T[6:0] ? 32'h0 : _GEN_119; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_121 = 7'h79 == _io_instruction_T[6:0] ? 32'h0 : _GEN_120; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_122 = 7'h7a == _io_instruction_T[6:0] ? 32'h0 : _GEN_121; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_123 = 7'h7b == _io_instruction_T[6:0] ? 32'h0 : _GEN_122; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_124 = 7'h7c == _io_instruction_T[6:0] ? 32'h0 : _GEN_123; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_125 = 7'h7d == _io_instruction_T[6:0] ? 32'h0 : _GEN_124; // @[instruction.scala 98:19 instruction.scala 98:19]
  wire [31:0] _GEN_126 = 7'h7e == _io_instruction_T[6:0] ? 32'h0 : _GEN_125; // @[instruction.scala 98:19 instruction.scala 98:19]
  assign io_instruction = reset ? 32'h0 : _GEN_126; // @[instruction.scala 19:23 instruction.scala 14:18 instruction.scala 98:19]
endmodule
module select(
  input  [7:0]  io_select_ctrl,
  input  [31:0] io_pc,
  input  [31:0] io_imm,
  input  [31:0] io_instruction,
  input  [31:0] io_data_read,
  input  [31:0] io_alu_out,
  input  [31:0] io_reg_read_data_1,
  input  [31:0] io_reg_read_data_2,
  output [31:0] io_data_addr,
  output [31:0] io_data_write,
  output [4:0]  io_reg_read_addr_1,
  output [4:0]  io_reg_read_addr_2,
  output [4:0]  io_reg_write_addr,
  output [31:0] io_reg_write_data,
  output [31:0] io_alu_src_1,
  output [31:0] io_alu_src_2,
  output [31:0] io_pc_imm
);
  wire  _T = 8'h7 == io_select_ctrl; // @[Conditional.scala 37:30]
  wire  _T_1 = 8'h1 == io_select_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _io_pc_imm_T_1 = io_pc + io_imm; // @[select.scala 50:28]
  wire [31:0] _io_pc_imm_T_3 = io_pc + 32'h4; // @[select.scala 53:28]
  wire [31:0] _GEN_0 = io_alu_out == 32'h1 ? _io_pc_imm_T_1 : _io_pc_imm_T_3; // @[select.scala 49:31 select.scala 50:19 select.scala 53:19]
  wire  _T_3 = 8'h0 == io_select_ctrl; // @[Conditional.scala 37:30]
  wire  _T_4 = 8'h4 == io_select_ctrl; // @[Conditional.scala 37:30]
  wire  _T_5 = 8'h2 == io_select_ctrl; // @[Conditional.scala 37:30]
  wire  _T_6 = 8'h3 == io_select_ctrl; // @[Conditional.scala 37:30]
  wire  _T_7 = 8'h8 == io_select_ctrl; // @[Conditional.scala 37:30]
  wire  _T_8 = 8'h5 == io_select_ctrl; // @[Conditional.scala 37:30]
  wire  _T_9 = 8'h6 == io_select_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_2 = _T_9 ? io_imm : io_reg_read_data_2; // @[Conditional.scala 39:67 select.scala 89:20 select.scala 36:16]
  wire [31:0] _GEN_3 = _T_9 ? io_alu_out : {{27'd0}, io_instruction[11:7]}; // @[Conditional.scala 39:67 select.scala 90:20 select.scala 29:17]
  wire [31:0] _GEN_4 = _T_9 ? io_reg_read_data_2 : io_alu_out; // @[Conditional.scala 39:67 select.scala 91:21 select.scala 30:17]
  wire [31:0] _GEN_6 = _T_8 ? io_reg_read_data_2 : _GEN_2; // @[Conditional.scala 39:67 select.scala 84:20]
  wire [31:0] _GEN_8 = _T_8 ? {{27'd0}, io_instruction[11:7]} : _GEN_3; // @[Conditional.scala 39:67 select.scala 29:17]
  wire [31:0] _GEN_9 = _T_8 ? io_alu_out : _GEN_4; // @[Conditional.scala 39:67 select.scala 30:17]
  wire [31:0] _GEN_10 = _T_7 ? io_imm : io_alu_out; // @[Conditional.scala 39:67 select.scala 80:25]
  wire [31:0] _GEN_12 = _T_7 ? io_reg_read_data_2 : _GEN_6; // @[Conditional.scala 39:67 select.scala 36:16]
  wire [31:0] _GEN_13 = _T_7 ? {{27'd0}, io_instruction[11:7]} : _GEN_8; // @[Conditional.scala 39:67 select.scala 29:17]
  wire [31:0] _GEN_14 = _T_7 ? io_alu_out : _GEN_9; // @[Conditional.scala 39:67 select.scala 30:17]
  wire [31:0] _GEN_16 = _T_6 ? io_imm : _GEN_12; // @[Conditional.scala 39:67 select.scala 75:20]
  wire [31:0] _GEN_17 = _T_6 ? io_alu_out : _GEN_13; // @[Conditional.scala 39:67 select.scala 76:20]
  wire [31:0] _GEN_18 = _T_6 ? io_data_read : _GEN_10; // @[Conditional.scala 39:67 select.scala 77:25]
  wire [31:0] _GEN_19 = _T_6 ? io_alu_out : _GEN_14; // @[Conditional.scala 39:67 select.scala 30:17]
  wire [31:0] _GEN_21 = _T_5 ? io_imm : _GEN_16; // @[Conditional.scala 39:67 select.scala 69:20]
  wire [31:0] _GEN_23 = _T_5 ? _io_pc_imm_T_3 : _GEN_18; // @[Conditional.scala 39:67 select.scala 71:25]
  wire [31:0] _GEN_24 = _T_5 ? {{27'd0}, io_instruction[11:7]} : _GEN_17; // @[Conditional.scala 39:67 select.scala 29:17]
  wire [31:0] _GEN_25 = _T_5 ? io_alu_out : _GEN_19; // @[Conditional.scala 39:67 select.scala 30:17]
  wire [31:0] _GEN_26 = _T_4 ? io_pc : io_reg_read_data_1; // @[Conditional.scala 39:67 select.scala 62:20]
  wire [31:0] _GEN_27 = _T_4 ? io_imm : _GEN_21; // @[Conditional.scala 39:67 select.scala 63:20]
  wire [31:0] _GEN_29 = _T_4 ? _io_pc_imm_T_3 : _GEN_23; // @[Conditional.scala 39:67 select.scala 65:25]
  wire [31:0] _GEN_30 = _T_4 ? {{27'd0}, io_instruction[11:7]} : _GEN_24; // @[Conditional.scala 39:67 select.scala 29:17]
  wire [31:0] _GEN_31 = _T_4 ? io_alu_out : _GEN_25; // @[Conditional.scala 39:67 select.scala 30:17]
  wire [31:0] _GEN_32 = _T_3 ? io_reg_read_data_1 : _GEN_26; // @[Conditional.scala 39:67 select.scala 57:20]
  wire [31:0] _GEN_33 = _T_3 ? io_imm : _GEN_27; // @[Conditional.scala 39:67 select.scala 58:20]
  wire [31:0] _GEN_34 = _T_3 ? io_alu_out : _GEN_31; // @[Conditional.scala 39:67 select.scala 59:21]
  wire [31:0] _GEN_36 = _T_3 ? io_alu_out : _GEN_29; // @[Conditional.scala 39:67 select.scala 34:21]
  wire [31:0] _GEN_37 = _T_3 ? {{27'd0}, io_instruction[11:7]} : _GEN_30; // @[Conditional.scala 39:67 select.scala 29:17]
  wire [31:0] _GEN_38 = _T_1 ? io_reg_read_data_1 : _GEN_32; // @[Conditional.scala 39:67 select.scala 47:20]
  wire [31:0] _GEN_39 = _T_1 ? io_reg_read_data_2 : _GEN_33; // @[Conditional.scala 39:67 select.scala 48:20]
  wire [31:0] _GEN_40 = _T_1 ? _GEN_0 : io_alu_out; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_41 = _T_1 ? io_alu_out : _GEN_34; // @[Conditional.scala 39:67 select.scala 30:17]
  wire [31:0] _GEN_42 = _T_1 ? io_alu_out : _GEN_36; // @[Conditional.scala 39:67 select.scala 34:21]
  wire [31:0] _GEN_43 = _T_1 ? {{27'd0}, io_instruction[11:7]} : _GEN_37; // @[Conditional.scala 39:67 select.scala 29:17]
  assign io_data_addr = _T ? {{27'd0}, io_instruction[11:7]} : _GEN_43; // @[Conditional.scala 40:58 select.scala 29:17]
  assign io_data_write = _T ? io_alu_out : _GEN_41; // @[Conditional.scala 40:58 select.scala 30:17]
  assign io_reg_read_addr_1 = io_instruction[19:15]; // @[select.scala 31:39]
  assign io_reg_read_addr_2 = io_instruction[24:20]; // @[select.scala 32:39]
  assign io_reg_write_addr = io_instruction[11:7]; // @[select.scala 33:38]
  assign io_reg_write_data = _T ? io_alu_out : _GEN_42; // @[Conditional.scala 40:58 select.scala 41:25]
  assign io_alu_src_1 = _T ? io_pc : _GEN_38; // @[Conditional.scala 40:58 select.scala 43:20]
  assign io_alu_src_2 = _T ? io_imm : _GEN_39; // @[Conditional.scala 40:58 select.scala 44:20]
  assign io_pc_imm = _T ? io_alu_out : _GEN_40; // @[Conditional.scala 40:58 select.scala 42:17]
endmodule
module reg_(
  input         clock,
  input         reset,
  input  [7:0]  io_reg_ctrl,
  input  [4:0]  io_reg_read_addr_1,
  input  [4:0]  io_reg_read_addr_2,
  input  [31:0] io_reg_write_data,
  input  [4:0]  io_reg_write_addr,
  output [31:0] io_reg_read_data_1,
  output [31:0] io_reg_read_data_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_1; // @[reg.scala 22:16]
  reg [31:0] reg_2; // @[reg.scala 22:16]
  reg [31:0] reg_3; // @[reg.scala 22:16]
  reg [31:0] reg_4; // @[reg.scala 22:16]
  reg [31:0] reg_5; // @[reg.scala 22:16]
  reg [31:0] reg_6; // @[reg.scala 22:16]
  reg [31:0] reg_7; // @[reg.scala 22:16]
  reg [31:0] reg_8; // @[reg.scala 22:16]
  reg [31:0] reg_9; // @[reg.scala 22:16]
  reg [31:0] reg_10; // @[reg.scala 22:16]
  reg [31:0] reg_11; // @[reg.scala 22:16]
  reg [31:0] reg_12; // @[reg.scala 22:16]
  reg [31:0] reg_13; // @[reg.scala 22:16]
  reg [31:0] reg_14; // @[reg.scala 22:16]
  reg [31:0] reg_15; // @[reg.scala 22:16]
  reg [31:0] reg_16; // @[reg.scala 22:16]
  reg [31:0] reg_17; // @[reg.scala 22:16]
  reg [31:0] reg_18; // @[reg.scala 22:16]
  reg [31:0] reg_19; // @[reg.scala 22:16]
  reg [31:0] reg_20; // @[reg.scala 22:16]
  reg [31:0] reg_21; // @[reg.scala 22:16]
  reg [31:0] reg_22; // @[reg.scala 22:16]
  reg [31:0] reg_23; // @[reg.scala 22:16]
  reg [31:0] reg_24; // @[reg.scala 22:16]
  reg [31:0] reg_25; // @[reg.scala 22:16]
  reg [31:0] reg_26; // @[reg.scala 22:16]
  reg [31:0] reg_27; // @[reg.scala 22:16]
  reg [31:0] reg_28; // @[reg.scala 22:16]
  reg [31:0] reg_29; // @[reg.scala 22:16]
  reg [31:0] reg_30; // @[reg.scala 22:16]
  reg [31:0] reg_31; // @[reg.scala 22:16]
  wire [31:0] _GEN_1 = 5'h1 == io_reg_read_addr_1 ? reg_1 : 32'h0; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_2 = 5'h2 == io_reg_read_addr_1 ? reg_2 : _GEN_1; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_3 = 5'h3 == io_reg_read_addr_1 ? reg_3 : _GEN_2; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_4 = 5'h4 == io_reg_read_addr_1 ? reg_4 : _GEN_3; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_5 = 5'h5 == io_reg_read_addr_1 ? reg_5 : _GEN_4; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_6 = 5'h6 == io_reg_read_addr_1 ? reg_6 : _GEN_5; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_7 = 5'h7 == io_reg_read_addr_1 ? reg_7 : _GEN_6; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_8 = 5'h8 == io_reg_read_addr_1 ? reg_8 : _GEN_7; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_9 = 5'h9 == io_reg_read_addr_1 ? reg_9 : _GEN_8; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_10 = 5'ha == io_reg_read_addr_1 ? reg_10 : _GEN_9; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_11 = 5'hb == io_reg_read_addr_1 ? reg_11 : _GEN_10; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_12 = 5'hc == io_reg_read_addr_1 ? reg_12 : _GEN_11; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_13 = 5'hd == io_reg_read_addr_1 ? reg_13 : _GEN_12; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_14 = 5'he == io_reg_read_addr_1 ? reg_14 : _GEN_13; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_15 = 5'hf == io_reg_read_addr_1 ? reg_15 : _GEN_14; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_16 = 5'h10 == io_reg_read_addr_1 ? reg_16 : _GEN_15; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_17 = 5'h11 == io_reg_read_addr_1 ? reg_17 : _GEN_16; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_18 = 5'h12 == io_reg_read_addr_1 ? reg_18 : _GEN_17; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_19 = 5'h13 == io_reg_read_addr_1 ? reg_19 : _GEN_18; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_20 = 5'h14 == io_reg_read_addr_1 ? reg_20 : _GEN_19; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_21 = 5'h15 == io_reg_read_addr_1 ? reg_21 : _GEN_20; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_22 = 5'h16 == io_reg_read_addr_1 ? reg_22 : _GEN_21; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_23 = 5'h17 == io_reg_read_addr_1 ? reg_23 : _GEN_22; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_24 = 5'h18 == io_reg_read_addr_1 ? reg_24 : _GEN_23; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_25 = 5'h19 == io_reg_read_addr_1 ? reg_25 : _GEN_24; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_26 = 5'h1a == io_reg_read_addr_1 ? reg_26 : _GEN_25; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_27 = 5'h1b == io_reg_read_addr_1 ? reg_27 : _GEN_26; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_28 = 5'h1c == io_reg_read_addr_1 ? reg_28 : _GEN_27; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_29 = 5'h1d == io_reg_read_addr_1 ? reg_29 : _GEN_28; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_30 = 5'h1e == io_reg_read_addr_1 ? reg_30 : _GEN_29; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_31 = 5'h1f == io_reg_read_addr_1 ? reg_31 : _GEN_30; // @[reg.scala 24:22 reg.scala 24:22]
  wire [31:0] _GEN_33 = 5'h1 == io_reg_read_addr_2 ? reg_1 : 32'h0; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_34 = 5'h2 == io_reg_read_addr_2 ? reg_2 : _GEN_33; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_35 = 5'h3 == io_reg_read_addr_2 ? reg_3 : _GEN_34; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_36 = 5'h4 == io_reg_read_addr_2 ? reg_4 : _GEN_35; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_37 = 5'h5 == io_reg_read_addr_2 ? reg_5 : _GEN_36; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_38 = 5'h6 == io_reg_read_addr_2 ? reg_6 : _GEN_37; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_39 = 5'h7 == io_reg_read_addr_2 ? reg_7 : _GEN_38; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_40 = 5'h8 == io_reg_read_addr_2 ? reg_8 : _GEN_39; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_41 = 5'h9 == io_reg_read_addr_2 ? reg_9 : _GEN_40; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_42 = 5'ha == io_reg_read_addr_2 ? reg_10 : _GEN_41; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_43 = 5'hb == io_reg_read_addr_2 ? reg_11 : _GEN_42; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_44 = 5'hc == io_reg_read_addr_2 ? reg_12 : _GEN_43; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_45 = 5'hd == io_reg_read_addr_2 ? reg_13 : _GEN_44; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_46 = 5'he == io_reg_read_addr_2 ? reg_14 : _GEN_45; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_47 = 5'hf == io_reg_read_addr_2 ? reg_15 : _GEN_46; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_48 = 5'h10 == io_reg_read_addr_2 ? reg_16 : _GEN_47; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_49 = 5'h11 == io_reg_read_addr_2 ? reg_17 : _GEN_48; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_50 = 5'h12 == io_reg_read_addr_2 ? reg_18 : _GEN_49; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_51 = 5'h13 == io_reg_read_addr_2 ? reg_19 : _GEN_50; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_52 = 5'h14 == io_reg_read_addr_2 ? reg_20 : _GEN_51; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_53 = 5'h15 == io_reg_read_addr_2 ? reg_21 : _GEN_52; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_54 = 5'h16 == io_reg_read_addr_2 ? reg_22 : _GEN_53; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_55 = 5'h17 == io_reg_read_addr_2 ? reg_23 : _GEN_54; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_56 = 5'h18 == io_reg_read_addr_2 ? reg_24 : _GEN_55; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_57 = 5'h19 == io_reg_read_addr_2 ? reg_25 : _GEN_56; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_58 = 5'h1a == io_reg_read_addr_2 ? reg_26 : _GEN_57; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_59 = 5'h1b == io_reg_read_addr_2 ? reg_27 : _GEN_58; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_60 = 5'h1c == io_reg_read_addr_2 ? reg_28 : _GEN_59; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_61 = 5'h1d == io_reg_read_addr_2 ? reg_29 : _GEN_60; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_62 = 5'h1e == io_reg_read_addr_2 ? reg_30 : _GEN_61; // @[reg.scala 25:22 reg.scala 25:22]
  wire [31:0] _GEN_63 = 5'h1f == io_reg_read_addr_2 ? reg_31 : _GEN_62; // @[reg.scala 25:22 reg.scala 25:22]
  wire  _T_1 = 8'h7 == io_reg_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_65 = 5'h1 == io_reg_write_addr ? io_reg_write_data : reg_1; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_66 = 5'h2 == io_reg_write_addr ? io_reg_write_data : reg_2; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_67 = 5'h3 == io_reg_write_addr ? io_reg_write_data : reg_3; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_68 = 5'h4 == io_reg_write_addr ? io_reg_write_data : reg_4; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_69 = 5'h5 == io_reg_write_addr ? io_reg_write_data : reg_5; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_70 = 5'h6 == io_reg_write_addr ? io_reg_write_data : reg_6; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_71 = 5'h7 == io_reg_write_addr ? io_reg_write_data : reg_7; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_72 = 5'h8 == io_reg_write_addr ? io_reg_write_data : reg_8; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_73 = 5'h9 == io_reg_write_addr ? io_reg_write_data : reg_9; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_74 = 5'ha == io_reg_write_addr ? io_reg_write_data : reg_10; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_75 = 5'hb == io_reg_write_addr ? io_reg_write_data : reg_11; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_76 = 5'hc == io_reg_write_addr ? io_reg_write_data : reg_12; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_77 = 5'hd == io_reg_write_addr ? io_reg_write_data : reg_13; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_78 = 5'he == io_reg_write_addr ? io_reg_write_data : reg_14; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_79 = 5'hf == io_reg_write_addr ? io_reg_write_data : reg_15; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_80 = 5'h10 == io_reg_write_addr ? io_reg_write_data : reg_16; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_81 = 5'h11 == io_reg_write_addr ? io_reg_write_data : reg_17; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_82 = 5'h12 == io_reg_write_addr ? io_reg_write_data : reg_18; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_83 = 5'h13 == io_reg_write_addr ? io_reg_write_data : reg_19; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_84 = 5'h14 == io_reg_write_addr ? io_reg_write_data : reg_20; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_85 = 5'h15 == io_reg_write_addr ? io_reg_write_data : reg_21; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_86 = 5'h16 == io_reg_write_addr ? io_reg_write_data : reg_22; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_87 = 5'h17 == io_reg_write_addr ? io_reg_write_data : reg_23; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_88 = 5'h18 == io_reg_write_addr ? io_reg_write_data : reg_24; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_89 = 5'h19 == io_reg_write_addr ? io_reg_write_data : reg_25; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_90 = 5'h1a == io_reg_write_addr ? io_reg_write_data : reg_26; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_91 = 5'h1b == io_reg_write_addr ? io_reg_write_data : reg_27; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_92 = 5'h1c == io_reg_write_addr ? io_reg_write_data : reg_28; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_93 = 5'h1d == io_reg_write_addr ? io_reg_write_data : reg_29; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_94 = 5'h1e == io_reg_write_addr ? io_reg_write_data : reg_30; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire [31:0] _GEN_95 = 5'h1f == io_reg_write_addr ? io_reg_write_data : reg_31; // @[reg.scala 34:30 reg.scala 34:30 reg.scala 22:16]
  wire  _T_2 = 8'h1 == io_reg_ctrl; // @[Conditional.scala 37:30]
  wire  _T_3 = 8'h0 == io_reg_ctrl; // @[Conditional.scala 37:30]
  wire  _T_4 = 8'h4 == io_reg_ctrl; // @[Conditional.scala 37:30]
  wire  _T_5 = 8'h2 == io_reg_ctrl; // @[Conditional.scala 37:30]
  wire  _T_6 = 8'h3 == io_reg_ctrl; // @[Conditional.scala 37:30]
  wire  _T_7 = 8'h8 == io_reg_ctrl; // @[Conditional.scala 37:30]
  wire  _T_8 = 8'h5 == io_reg_ctrl; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_290 = _T_8 ? _GEN_65 : reg_1; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_291 = _T_8 ? _GEN_66 : reg_2; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_292 = _T_8 ? _GEN_67 : reg_3; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_293 = _T_8 ? _GEN_68 : reg_4; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_294 = _T_8 ? _GEN_69 : reg_5; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_295 = _T_8 ? _GEN_70 : reg_6; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_296 = _T_8 ? _GEN_71 : reg_7; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_297 = _T_8 ? _GEN_72 : reg_8; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_298 = _T_8 ? _GEN_73 : reg_9; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_299 = _T_8 ? _GEN_74 : reg_10; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_300 = _T_8 ? _GEN_75 : reg_11; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_301 = _T_8 ? _GEN_76 : reg_12; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_302 = _T_8 ? _GEN_77 : reg_13; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_303 = _T_8 ? _GEN_78 : reg_14; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_304 = _T_8 ? _GEN_79 : reg_15; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_305 = _T_8 ? _GEN_80 : reg_16; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_306 = _T_8 ? _GEN_81 : reg_17; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_307 = _T_8 ? _GEN_82 : reg_18; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_308 = _T_8 ? _GEN_83 : reg_19; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_309 = _T_8 ? _GEN_84 : reg_20; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_310 = _T_8 ? _GEN_85 : reg_21; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_311 = _T_8 ? _GEN_86 : reg_22; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_312 = _T_8 ? _GEN_87 : reg_23; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_313 = _T_8 ? _GEN_88 : reg_24; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_314 = _T_8 ? _GEN_89 : reg_25; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_315 = _T_8 ? _GEN_90 : reg_26; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_316 = _T_8 ? _GEN_91 : reg_27; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_317 = _T_8 ? _GEN_92 : reg_28; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_318 = _T_8 ? _GEN_93 : reg_29; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_319 = _T_8 ? _GEN_94 : reg_30; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_320 = _T_8 ? _GEN_95 : reg_31; // @[Conditional.scala 39:67 reg.scala 22:16]
  wire [31:0] _GEN_322 = _T_7 ? _GEN_65 : _GEN_290; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_323 = _T_7 ? _GEN_66 : _GEN_291; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_324 = _T_7 ? _GEN_67 : _GEN_292; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_325 = _T_7 ? _GEN_68 : _GEN_293; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_326 = _T_7 ? _GEN_69 : _GEN_294; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_327 = _T_7 ? _GEN_70 : _GEN_295; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_328 = _T_7 ? _GEN_71 : _GEN_296; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_329 = _T_7 ? _GEN_72 : _GEN_297; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_330 = _T_7 ? _GEN_73 : _GEN_298; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_331 = _T_7 ? _GEN_74 : _GEN_299; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_332 = _T_7 ? _GEN_75 : _GEN_300; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_333 = _T_7 ? _GEN_76 : _GEN_301; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_334 = _T_7 ? _GEN_77 : _GEN_302; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_335 = _T_7 ? _GEN_78 : _GEN_303; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_336 = _T_7 ? _GEN_79 : _GEN_304; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_337 = _T_7 ? _GEN_80 : _GEN_305; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_338 = _T_7 ? _GEN_81 : _GEN_306; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_339 = _T_7 ? _GEN_82 : _GEN_307; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_340 = _T_7 ? _GEN_83 : _GEN_308; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_341 = _T_7 ? _GEN_84 : _GEN_309; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_342 = _T_7 ? _GEN_85 : _GEN_310; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_343 = _T_7 ? _GEN_86 : _GEN_311; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_344 = _T_7 ? _GEN_87 : _GEN_312; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_345 = _T_7 ? _GEN_88 : _GEN_313; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_346 = _T_7 ? _GEN_89 : _GEN_314; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_347 = _T_7 ? _GEN_90 : _GEN_315; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_348 = _T_7 ? _GEN_91 : _GEN_316; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_349 = _T_7 ? _GEN_92 : _GEN_317; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_350 = _T_7 ? _GEN_93 : _GEN_318; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_351 = _T_7 ? _GEN_94 : _GEN_319; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_352 = _T_7 ? _GEN_95 : _GEN_320; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_354 = _T_6 ? _GEN_65 : _GEN_322; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_355 = _T_6 ? _GEN_66 : _GEN_323; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_356 = _T_6 ? _GEN_67 : _GEN_324; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_357 = _T_6 ? _GEN_68 : _GEN_325; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_358 = _T_6 ? _GEN_69 : _GEN_326; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_359 = _T_6 ? _GEN_70 : _GEN_327; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_360 = _T_6 ? _GEN_71 : _GEN_328; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_361 = _T_6 ? _GEN_72 : _GEN_329; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_362 = _T_6 ? _GEN_73 : _GEN_330; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_363 = _T_6 ? _GEN_74 : _GEN_331; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_364 = _T_6 ? _GEN_75 : _GEN_332; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_365 = _T_6 ? _GEN_76 : _GEN_333; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_366 = _T_6 ? _GEN_77 : _GEN_334; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_367 = _T_6 ? _GEN_78 : _GEN_335; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_368 = _T_6 ? _GEN_79 : _GEN_336; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_369 = _T_6 ? _GEN_80 : _GEN_337; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_370 = _T_6 ? _GEN_81 : _GEN_338; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_371 = _T_6 ? _GEN_82 : _GEN_339; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_372 = _T_6 ? _GEN_83 : _GEN_340; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_373 = _T_6 ? _GEN_84 : _GEN_341; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_374 = _T_6 ? _GEN_85 : _GEN_342; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_375 = _T_6 ? _GEN_86 : _GEN_343; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_376 = _T_6 ? _GEN_87 : _GEN_344; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_377 = _T_6 ? _GEN_88 : _GEN_345; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_378 = _T_6 ? _GEN_89 : _GEN_346; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_379 = _T_6 ? _GEN_90 : _GEN_347; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_380 = _T_6 ? _GEN_91 : _GEN_348; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_381 = _T_6 ? _GEN_92 : _GEN_349; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_382 = _T_6 ? _GEN_93 : _GEN_350; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_383 = _T_6 ? _GEN_94 : _GEN_351; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_384 = _T_6 ? _GEN_95 : _GEN_352; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_386 = _T_5 ? _GEN_65 : _GEN_354; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_387 = _T_5 ? _GEN_66 : _GEN_355; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_388 = _T_5 ? _GEN_67 : _GEN_356; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_389 = _T_5 ? _GEN_68 : _GEN_357; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_390 = _T_5 ? _GEN_69 : _GEN_358; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_391 = _T_5 ? _GEN_70 : _GEN_359; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_392 = _T_5 ? _GEN_71 : _GEN_360; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_393 = _T_5 ? _GEN_72 : _GEN_361; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_394 = _T_5 ? _GEN_73 : _GEN_362; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_395 = _T_5 ? _GEN_74 : _GEN_363; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_396 = _T_5 ? _GEN_75 : _GEN_364; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_397 = _T_5 ? _GEN_76 : _GEN_365; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_398 = _T_5 ? _GEN_77 : _GEN_366; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_399 = _T_5 ? _GEN_78 : _GEN_367; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_400 = _T_5 ? _GEN_79 : _GEN_368; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_401 = _T_5 ? _GEN_80 : _GEN_369; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_402 = _T_5 ? _GEN_81 : _GEN_370; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_403 = _T_5 ? _GEN_82 : _GEN_371; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_404 = _T_5 ? _GEN_83 : _GEN_372; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_405 = _T_5 ? _GEN_84 : _GEN_373; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_406 = _T_5 ? _GEN_85 : _GEN_374; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_407 = _T_5 ? _GEN_86 : _GEN_375; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_408 = _T_5 ? _GEN_87 : _GEN_376; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_409 = _T_5 ? _GEN_88 : _GEN_377; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_410 = _T_5 ? _GEN_89 : _GEN_378; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_411 = _T_5 ? _GEN_90 : _GEN_379; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_412 = _T_5 ? _GEN_91 : _GEN_380; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_413 = _T_5 ? _GEN_92 : _GEN_381; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_414 = _T_5 ? _GEN_93 : _GEN_382; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_415 = _T_5 ? _GEN_94 : _GEN_383; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_416 = _T_5 ? _GEN_95 : _GEN_384; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_418 = _T_4 ? _GEN_65 : _GEN_386; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_419 = _T_4 ? _GEN_66 : _GEN_387; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_420 = _T_4 ? _GEN_67 : _GEN_388; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_421 = _T_4 ? _GEN_68 : _GEN_389; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_422 = _T_4 ? _GEN_69 : _GEN_390; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_423 = _T_4 ? _GEN_70 : _GEN_391; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_424 = _T_4 ? _GEN_71 : _GEN_392; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_425 = _T_4 ? _GEN_72 : _GEN_393; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_426 = _T_4 ? _GEN_73 : _GEN_394; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_427 = _T_4 ? _GEN_74 : _GEN_395; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_428 = _T_4 ? _GEN_75 : _GEN_396; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_429 = _T_4 ? _GEN_76 : _GEN_397; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_430 = _T_4 ? _GEN_77 : _GEN_398; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_431 = _T_4 ? _GEN_78 : _GEN_399; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_432 = _T_4 ? _GEN_79 : _GEN_400; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_433 = _T_4 ? _GEN_80 : _GEN_401; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_434 = _T_4 ? _GEN_81 : _GEN_402; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_435 = _T_4 ? _GEN_82 : _GEN_403; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_436 = _T_4 ? _GEN_83 : _GEN_404; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_437 = _T_4 ? _GEN_84 : _GEN_405; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_438 = _T_4 ? _GEN_85 : _GEN_406; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_439 = _T_4 ? _GEN_86 : _GEN_407; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_440 = _T_4 ? _GEN_87 : _GEN_408; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_441 = _T_4 ? _GEN_88 : _GEN_409; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_442 = _T_4 ? _GEN_89 : _GEN_410; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_443 = _T_4 ? _GEN_90 : _GEN_411; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_444 = _T_4 ? _GEN_91 : _GEN_412; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_445 = _T_4 ? _GEN_92 : _GEN_413; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_446 = _T_4 ? _GEN_93 : _GEN_414; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_447 = _T_4 ? _GEN_94 : _GEN_415; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_448 = _T_4 ? _GEN_95 : _GEN_416; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_545 = io_reg_read_addr_1 == 5'h0 ? 32'h0 : _GEN_31; // @[reg.scala 70:35 reg.scala 71:24 reg.scala 24:22]
  wire [31:0] _GEN_546 = io_reg_read_addr_2 == 5'h0 ? 32'h0 : _GEN_63; // @[reg.scala 73:35 reg.scala 74:24 reg.scala 25:22]
  assign io_reg_read_data_1 = reset ? _GEN_31 : _GEN_545; // @[reg.scala 27:23 reg.scala 24:22]
  assign io_reg_read_data_2 = reset ? _GEN_63 : _GEN_546; // @[reg.scala 27:23 reg.scala 25:22]
  always @(posedge clock) begin
    if (reset) begin // @[reg.scala 27:23]
      reg_1 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_1 <= _GEN_65;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_1 <= _GEN_65;
      end else begin
        reg_1 <= _GEN_418;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_2 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_2 <= _GEN_66;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_2 <= _GEN_66;
      end else begin
        reg_2 <= _GEN_419;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_3 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_3 <= _GEN_67;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_3 <= _GEN_67;
      end else begin
        reg_3 <= _GEN_420;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_4 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_4 <= _GEN_68;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_4 <= _GEN_68;
      end else begin
        reg_4 <= _GEN_421;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_5 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_5 <= _GEN_69;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_5 <= _GEN_69;
      end else begin
        reg_5 <= _GEN_422;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_6 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_6 <= _GEN_70;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_6 <= _GEN_70;
      end else begin
        reg_6 <= _GEN_423;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_7 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_7 <= _GEN_71;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_7 <= _GEN_71;
      end else begin
        reg_7 <= _GEN_424;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_8 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_8 <= _GEN_72;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_8 <= _GEN_72;
      end else begin
        reg_8 <= _GEN_425;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_9 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_9 <= _GEN_73;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_9 <= _GEN_73;
      end else begin
        reg_9 <= _GEN_426;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_10 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_10 <= _GEN_74;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_10 <= _GEN_74;
      end else begin
        reg_10 <= _GEN_427;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_11 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_11 <= _GEN_75;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_11 <= _GEN_75;
      end else begin
        reg_11 <= _GEN_428;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_12 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_12 <= _GEN_76;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_12 <= _GEN_76;
      end else begin
        reg_12 <= _GEN_429;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_13 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_13 <= _GEN_77;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_13 <= _GEN_77;
      end else begin
        reg_13 <= _GEN_430;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_14 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_14 <= _GEN_78;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_14 <= _GEN_78;
      end else begin
        reg_14 <= _GEN_431;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_15 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_15 <= _GEN_79;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_15 <= _GEN_79;
      end else begin
        reg_15 <= _GEN_432;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_16 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_16 <= _GEN_80;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_16 <= _GEN_80;
      end else begin
        reg_16 <= _GEN_433;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_17 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_17 <= _GEN_81;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_17 <= _GEN_81;
      end else begin
        reg_17 <= _GEN_434;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_18 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_18 <= _GEN_82;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_18 <= _GEN_82;
      end else begin
        reg_18 <= _GEN_435;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_19 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_19 <= _GEN_83;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_19 <= _GEN_83;
      end else begin
        reg_19 <= _GEN_436;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_20 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_20 <= _GEN_84;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_20 <= _GEN_84;
      end else begin
        reg_20 <= _GEN_437;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_21 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_21 <= _GEN_85;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_21 <= _GEN_85;
      end else begin
        reg_21 <= _GEN_438;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_22 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_22 <= _GEN_86;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_22 <= _GEN_86;
      end else begin
        reg_22 <= _GEN_439;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_23 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_23 <= _GEN_87;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_23 <= _GEN_87;
      end else begin
        reg_23 <= _GEN_440;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_24 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_24 <= _GEN_88;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_24 <= _GEN_88;
      end else begin
        reg_24 <= _GEN_441;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_25 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_25 <= _GEN_89;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_25 <= _GEN_89;
      end else begin
        reg_25 <= _GEN_442;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_26 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_26 <= _GEN_90;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_26 <= _GEN_90;
      end else begin
        reg_26 <= _GEN_443;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_27 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_27 <= _GEN_91;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_27 <= _GEN_91;
      end else begin
        reg_27 <= _GEN_444;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_28 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_28 <= _GEN_92;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_28 <= _GEN_92;
      end else begin
        reg_28 <= _GEN_445;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_29 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_29 <= _GEN_93;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_29 <= _GEN_93;
      end else begin
        reg_29 <= _GEN_446;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_30 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_30 <= _GEN_94;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_30 <= _GEN_94;
      end else begin
        reg_30 <= _GEN_447;
      end
    end
    if (reset) begin // @[reg.scala 27:23]
      reg_31 <= 32'h0; // @[reg.scala 29:16]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      reg_31 <= _GEN_95;
    end else if (!(_T_2)) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Conditional.scala 39:67]
        reg_31 <= _GEN_95;
      end else begin
        reg_31 <= _GEN_448;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_1 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_2 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_3 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_7 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_8 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_9 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_10 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_11 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_12 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_13 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_14 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_15 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_16 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_17 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_18 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_19 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_20 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_21 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_22 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_23 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_24 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_25 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_26 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_27 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_28 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_29 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_30 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_31 = _RAND_30[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CPU(
  input         clock,
  input         reset,
  output [31:0] io_out
);
  wire  mod_pc_clock; // @[cpu.scala 37:22]
  wire  mod_pc_reset; // @[cpu.scala 37:22]
  wire [7:0] mod_pc_io_pc_ctrl; // @[cpu.scala 37:22]
  wire [31:0] mod_pc_io_pc_imm; // @[cpu.scala 37:22]
  wire [31:0] mod_pc_io_pc; // @[cpu.scala 37:22]
  wire [7:0] mod_alu_io_alu_ctrl; // @[cpu.scala 41:23]
  wire [31:0] mod_alu_io_alu_src_1; // @[cpu.scala 41:23]
  wire [31:0] mod_alu_io_alu_src_2; // @[cpu.scala 41:23]
  wire [31:0] mod_alu_io_alu_out; // @[cpu.scala 41:23]
  wire [31:0] mod_ctrl_io_instruction; // @[cpu.scala 46:24]
  wire [7:0] mod_ctrl_io_pc_ctrl; // @[cpu.scala 46:24]
  wire [7:0] mod_ctrl_io_imm_ctrl; // @[cpu.scala 46:24]
  wire [7:0] mod_ctrl_io_data_ctrl; // @[cpu.scala 46:24]
  wire [7:0] mod_ctrl_io_select_ctrl; // @[cpu.scala 46:24]
  wire [7:0] mod_ctrl_io_reg_ctrl; // @[cpu.scala 46:24]
  wire [7:0] mod_ctrl_io_alu_ctrl; // @[cpu.scala 46:24]
  wire  mod_data_clock; // @[cpu.scala 54:24]
  wire  mod_data_reset; // @[cpu.scala 54:24]
  wire [7:0] mod_data_io_data_ctrl; // @[cpu.scala 54:24]
  wire [31:0] mod_data_io_data_addr; // @[cpu.scala 54:24]
  wire [31:0] mod_data_io_data_write; // @[cpu.scala 54:24]
  wire [31:0] mod_data_io_data_read; // @[cpu.scala 54:24]
  wire [7:0] mod_imm_gen_io_imm_ctrl; // @[cpu.scala 59:27]
  wire [31:0] mod_imm_gen_io_instruction; // @[cpu.scala 59:27]
  wire [31:0] mod_imm_gen_io_imm; // @[cpu.scala 59:27]
  wire  mod_instruction_reset; // @[cpu.scala 63:31]
  wire [31:0] mod_instruction_io_pc; // @[cpu.scala 63:31]
  wire [31:0] mod_instruction_io_instruction; // @[cpu.scala 63:31]
  wire [7:0] mod_select_io_select_ctrl; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_pc; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_imm; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_instruction; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_data_read; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_alu_out; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_reg_read_data_1; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_reg_read_data_2; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_data_addr; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_data_write; // @[cpu.scala 66:26]
  wire [4:0] mod_select_io_reg_read_addr_1; // @[cpu.scala 66:26]
  wire [4:0] mod_select_io_reg_read_addr_2; // @[cpu.scala 66:26]
  wire [4:0] mod_select_io_reg_write_addr; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_reg_write_data; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_alu_src_1; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_alu_src_2; // @[cpu.scala 66:26]
  wire [31:0] mod_select_io_pc_imm; // @[cpu.scala 66:26]
  wire  mod_reg_clock; // @[cpu.scala 84:23]
  wire  mod_reg_reset; // @[cpu.scala 84:23]
  wire [7:0] mod_reg_io_reg_ctrl; // @[cpu.scala 84:23]
  wire [4:0] mod_reg_io_reg_read_addr_1; // @[cpu.scala 84:23]
  wire [4:0] mod_reg_io_reg_read_addr_2; // @[cpu.scala 84:23]
  wire [31:0] mod_reg_io_reg_write_data; // @[cpu.scala 84:23]
  wire [4:0] mod_reg_io_reg_write_addr; // @[cpu.scala 84:23]
  wire [31:0] mod_reg_io_reg_read_data_1; // @[cpu.scala 84:23]
  wire [31:0] mod_reg_io_reg_read_data_2; // @[cpu.scala 84:23]
  wire [4:0] data_addr = mod_select_io_data_addr[4:0]; // @[cpu.scala 17:23 cpu.scala 75:15]
  pc mod_pc ( // @[cpu.scala 37:22]
    .clock(mod_pc_clock),
    .reset(mod_pc_reset),
    .io_pc_ctrl(mod_pc_io_pc_ctrl),
    .io_pc_imm(mod_pc_io_pc_imm),
    .io_pc(mod_pc_io_pc)
  );
  alu mod_alu ( // @[cpu.scala 41:23]
    .io_alu_ctrl(mod_alu_io_alu_ctrl),
    .io_alu_src_1(mod_alu_io_alu_src_1),
    .io_alu_src_2(mod_alu_io_alu_src_2),
    .io_alu_out(mod_alu_io_alu_out)
  );
  ctrl mod_ctrl ( // @[cpu.scala 46:24]
    .io_instruction(mod_ctrl_io_instruction),
    .io_pc_ctrl(mod_ctrl_io_pc_ctrl),
    .io_imm_ctrl(mod_ctrl_io_imm_ctrl),
    .io_data_ctrl(mod_ctrl_io_data_ctrl),
    .io_select_ctrl(mod_ctrl_io_select_ctrl),
    .io_reg_ctrl(mod_ctrl_io_reg_ctrl),
    .io_alu_ctrl(mod_ctrl_io_alu_ctrl)
  );
  data mod_data ( // @[cpu.scala 54:24]
    .clock(mod_data_clock),
    .reset(mod_data_reset),
    .io_data_ctrl(mod_data_io_data_ctrl),
    .io_data_addr(mod_data_io_data_addr),
    .io_data_write(mod_data_io_data_write),
    .io_data_read(mod_data_io_data_read)
  );
  imm_gen mod_imm_gen ( // @[cpu.scala 59:27]
    .io_imm_ctrl(mod_imm_gen_io_imm_ctrl),
    .io_instruction(mod_imm_gen_io_instruction),
    .io_imm(mod_imm_gen_io_imm)
  );
  instruction mod_instruction ( // @[cpu.scala 63:31]
    .reset(mod_instruction_reset),
    .io_pc(mod_instruction_io_pc),
    .io_instruction(mod_instruction_io_instruction)
  );
  select mod_select ( // @[cpu.scala 66:26]
    .io_select_ctrl(mod_select_io_select_ctrl),
    .io_pc(mod_select_io_pc),
    .io_imm(mod_select_io_imm),
    .io_instruction(mod_select_io_instruction),
    .io_data_read(mod_select_io_data_read),
    .io_alu_out(mod_select_io_alu_out),
    .io_reg_read_data_1(mod_select_io_reg_read_data_1),
    .io_reg_read_data_2(mod_select_io_reg_read_data_2),
    .io_data_addr(mod_select_io_data_addr),
    .io_data_write(mod_select_io_data_write),
    .io_reg_read_addr_1(mod_select_io_reg_read_addr_1),
    .io_reg_read_addr_2(mod_select_io_reg_read_addr_2),
    .io_reg_write_addr(mod_select_io_reg_write_addr),
    .io_reg_write_data(mod_select_io_reg_write_data),
    .io_alu_src_1(mod_select_io_alu_src_1),
    .io_alu_src_2(mod_select_io_alu_src_2),
    .io_pc_imm(mod_select_io_pc_imm)
  );
  reg_ mod_reg ( // @[cpu.scala 84:23]
    .clock(mod_reg_clock),
    .reset(mod_reg_reset),
    .io_reg_ctrl(mod_reg_io_reg_ctrl),
    .io_reg_read_addr_1(mod_reg_io_reg_read_addr_1),
    .io_reg_read_addr_2(mod_reg_io_reg_read_addr_2),
    .io_reg_write_data(mod_reg_io_reg_write_data),
    .io_reg_write_addr(mod_reg_io_reg_write_addr),
    .io_reg_read_data_1(mod_reg_io_reg_read_data_1),
    .io_reg_read_data_2(mod_reg_io_reg_read_data_2)
  );
  assign io_out = mod_instruction_io_instruction; // @[cpu.scala 93:10]
  assign mod_pc_clock = clock;
  assign mod_pc_reset = reset;
  assign mod_pc_io_pc_ctrl = mod_ctrl_io_pc_ctrl; // @[cpu.scala 26:21 cpu.scala 48:13]
  assign mod_pc_io_pc_imm = mod_select_io_pc_imm; // @[cpu.scala 25:20 cpu.scala 83:12]
  assign mod_alu_io_alu_ctrl = mod_ctrl_io_alu_ctrl; // @[cpu.scala 31:22 cpu.scala 53:14]
  assign mod_alu_io_alu_src_1 = mod_select_io_alu_src_1; // @[cpu.scala 23:23 cpu.scala 81:15]
  assign mod_alu_io_alu_src_2 = mod_select_io_alu_src_2; // @[cpu.scala 24:23 cpu.scala 82:15]
  assign mod_ctrl_io_instruction = mod_instruction_io_instruction; // @[cpu.scala 14:25 cpu.scala 65:17]
  assign mod_data_clock = clock;
  assign mod_data_reset = reset;
  assign mod_data_io_data_ctrl = mod_ctrl_io_data_ctrl; // @[cpu.scala 28:23 cpu.scala 50:15]
  assign mod_data_io_data_addr = {{27'd0}, data_addr}; // @[cpu.scala 17:23 cpu.scala 75:15]
  assign mod_data_io_data_write = mod_select_io_data_write; // @[cpu.scala 18:24 cpu.scala 76:16]
  assign mod_imm_gen_io_imm_ctrl = mod_ctrl_io_imm_ctrl; // @[cpu.scala 27:22 cpu.scala 49:14]
  assign mod_imm_gen_io_instruction = mod_instruction_io_instruction; // @[cpu.scala 14:25 cpu.scala 65:17]
  assign mod_instruction_reset = reset;
  assign mod_instruction_io_pc = mod_pc_io_pc; // @[cpu.scala 13:16 cpu.scala 40:8]
  assign mod_select_io_select_ctrl = mod_ctrl_io_select_ctrl; // @[cpu.scala 29:25 cpu.scala 51:17]
  assign mod_select_io_pc = mod_pc_io_pc; // @[cpu.scala 13:16 cpu.scala 40:8]
  assign mod_select_io_imm = mod_imm_gen_io_imm; // @[cpu.scala 15:17 cpu.scala 62:9]
  assign mod_select_io_instruction = mod_instruction_io_instruction; // @[cpu.scala 14:25 cpu.scala 65:17]
  assign mod_select_io_data_read = mod_data_io_data_read; // @[cpu.scala 16:23 cpu.scala 58:15]
  assign mod_select_io_alu_out = mod_alu_io_alu_out; // @[cpu.scala 34:21 cpu.scala 45:13]
  assign mod_select_io_reg_read_data_1 = mod_reg_io_reg_read_data_1; // @[cpu.scala 32:29 cpu.scala 90:21]
  assign mod_select_io_reg_read_data_2 = mod_reg_io_reg_read_data_2; // @[cpu.scala 33:29 cpu.scala 91:21]
  assign mod_reg_clock = clock;
  assign mod_reg_reset = reset;
  assign mod_reg_io_reg_ctrl = mod_ctrl_io_reg_ctrl; // @[cpu.scala 30:22 cpu.scala 52:14]
  assign mod_reg_io_reg_read_addr_1 = mod_select_io_reg_read_addr_1; // @[cpu.scala 19:29 cpu.scala 77:21]
  assign mod_reg_io_reg_read_addr_2 = mod_select_io_reg_read_addr_2; // @[cpu.scala 20:29 cpu.scala 78:21]
  assign mod_reg_io_reg_write_data = mod_select_io_reg_write_data; // @[cpu.scala 22:28 cpu.scala 80:20]
  assign mod_reg_io_reg_write_addr = mod_select_io_reg_write_addr; // @[cpu.scala 21:28 cpu.scala 79:20]
endmodule
